library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is
    generic(
        AddrWidth   : integer := 13
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end monitor;

architecture rtl of monitor is
    type rom8192x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom8192x8 := (
         x"31",  x"c0",  x"eb",  x"21",  x"54",  x"00",  x"11",  x"00", -- 0000
         x"80",  x"cd",  x"0f",  x"00",  x"c3",  x"10",  x"80",  x"3e", -- 0008
         x"80",  x"ed",  x"a0",  x"cd",  x"4e",  x"00",  x"30",  x"f9", -- 0010
         x"d5",  x"01",  x"00",  x"00",  x"50",  x"14",  x"cd",  x"4e", -- 0018
         x"00",  x"30",  x"fa",  x"d4",  x"4e",  x"00",  x"cb",  x"11", -- 0020
         x"cb",  x"10",  x"38",  x"1f",  x"15",  x"20",  x"f4",  x"03", -- 0028
         x"5e",  x"23",  x"cb",  x"33",  x"30",  x"0c",  x"16",  x"10", -- 0030
         x"cd",  x"4e",  x"00",  x"cb",  x"12",  x"30",  x"f9",  x"14", -- 0038
         x"cb",  x"3a",  x"cb",  x"1b",  x"e3",  x"e5",  x"ed",  x"52", -- 0040
         x"d1",  x"ed",  x"b0",  x"e1",  x"30",  x"c5",  x"87",  x"c0", -- 0048
         x"7e",  x"23",  x"17",  x"c9",  x"c3",  x"04",  x"0c",  x"80", -- 0050
         x"53",  x"44",  x"20",  x"80",  x"00",  x"00",  x"3e",  x"01", -- 0058
         x"d3",  x"02",  x"00",  x"31",  x"00",  x"c0",  x"cd",  x"0c", -- 0060
         x"af",  x"cd",  x"2a",  x"07",  x"87",  x"c3",  x"03",  x"f0", -- 0068
         x"00",  x"00",  x"80",  x"13",  x"02",  x"cf",  x"c9",  x"3e", -- 0070
         x"00",  x"cf",  x"76",  x"03",  x"18",  x"fd",  x"dd",  x"e5", -- 0078
         x"dd",  x"21",  x"0f",  x"00",  x"dd",  x"39",  x"f5",  x"dd", -- 0080
         x"7e",  x"04",  x"dd",  x"77",  x"6c",  x"fe",  x"05",  x"05", -- 0088
         x"05",  x"ff",  x"e1",  x"00",  x"e5",  x"56",  x"23",  x"66", -- 0090
         x"dd",  x"4e",  x"06",  x"06",  x"00",  x"00",  x"7a",  x"a9", -- 0098
         x"5f",  x"7c",  x"a8",  x"57",  x"26",  x"00",  x"00",  x"cb", -- 00A0
         x"7c",  x"28",  x"19",  x"6b",  x"42",  x"cb",  x"00",  x"28", -- 00A8
         x"cb",  x"1d",  x"cb",  x"43",  x"28",  x"0a",  x"7d",  x"00", -- 00B0
         x"ee",  x"01",  x"5f",  x"78",  x"ee",  x"a0",  x"57",  x"18", -- 00B8
         x"03",  x"02",  x"5d",  x"50",  x"24",  x"18",  x"e3",  x"2e", -- 00C0
         x"00",  x"73",  x"23",  x"72",  x"f1",  x"dd",  x"e1",  x"c9", -- 00C8
         x"f5",  x"00",  x"21",  x"04",  x"00",  x"39",  x"4e",  x"23", -- 00D0
         x"46",  x"c5",  x"00",  x"cd",  x"81",  x"a2",  x"f1",  x"55", -- 00D8
         x"7a",  x"b7",  x"20",  x"78",  x"3e",  x"5b",  x"10",  x"e5", -- 00E0
         x"21",  x"0a",  x"96",  x"15",  x"70",  x"07",  x"cd",  x"78", -- 00E8
         x"a3",  x"f1",  x"d6",  x"00",  x"55",  x"1b",  x"7e",  x"00", -- 00F0
         x"fd",  x"21",  x"08",  x"00",  x"fd",  x"39",  x"fd",  x"96", -- 00F8
         x"04",  x"00",  x"20",  x"10",  x"21",  x"01",  x"50",  x"0f", -- 0100
         x"01",  x"28",  x"02",  x"04",  x"16",  x"01",  x"6a",  x"f1", -- 0108
         x"c9",  x"40",  x"9f",  x"60",  x"00",  x"21",  x"26",  x"b2", -- 0110
         x"36",  x"00",  x"2d",  x"21",  x"27",  x"04",  x"2a",  x"6b", -- 0118
         x"04",  x"2b",  x"04",  x"5a",  x"28",  x"04",  x"29",  x"d6", -- 0120
         x"04",  x"15",  x"04",  x"1e",  x"f6",  x"04",  x"2c",  x"6e", -- 0128
         x"c9",  x"02",  x"66",  x"05",  x"e5",  x"c0",  x"83",  x"dd", -- 0130
         x"75",  x"02",  x"fc",  x"7d",  x"b7",  x"c2",  x"64",  x"84", -- 0138
         x"fc",  x"6a",  x"0b",  x"dd",  x"00",  x"74",  x"ff",  x"eb", -- 0140
         x"21",  x"1a",  x"b1",  x"07",  x"d5",  x"01",  x"10",  x"00", -- 0148
         x"c5",  x"1f",  x"61",  x"85",  x"13",  x"21",  x"d8",  x"16", -- 0150
         x"15",  x"01",  x"85",  x"84",  x"a2",  x"19",  x"a6",  x"ac", -- 0158
         x"20",  x"19",  x"46",  x"83",  x"32",  x"dd",  x"5e",  x"37", -- 0160
         x"56",  x"ff",  x"44",  x"36",  x"81",  x"69",  x"36",  x"28", -- 0168
         x"0e",  x"88",  x"ae",  x"fa",  x"d6",  x"81",  x"31",  x"20", -- 0170
         x"07",  x"06",  x"fb",  x"b7",  x"ca",  x"bc",  x"29",  x"3a", -- 0178
         x"23",  x"bc",  x"40",  x"fd",  x"3d",  x"c2",  x"69",  x"82", -- 0180
         x"3a",  x"0b",  x"1b",  x"b1",  x"d6",  x"d3",  x"07",  x"4c", -- 0188
         x"1c",  x"07",  x"1d",  x"94",  x"07",  x"21",  x"96",  x"62", -- 0190
         x"84",  x"40",  x"c0",  x"8b",  x"f1",  x"c0",  x"a7",  x"01", -- 0198
         x"1e",  x"c2",  x"e8",  x"80",  x"b4",  x"d5",  x"16",  x"c2", -- 01A0
         x"06",  x"19",  x"d1",  x"4b",  x"0c",  x"ab",  x"00",  x"63", -- 01A8
         x"f1",  x"16",  x"09",  x"82",  x"20",  x"77",  x"00",  x"1c", -- 01B0
         x"7b",  x"d6",  x"15",  x"08",  x"38",  x"e1",  x"1d",  x"a4", -- 01B8
         x"1c",  x"19",  x"da",  x"0b",  x"35",  x"00",  x"26",  x"0a", -- 01C0
         x"e3",  x"33",  x"cd",  x"aa",  x"8b",  x"33",  x"b1",  x"87", -- 01C8
         x"58",  x"01",  x"87",  x"8b",  x"04",  x"21",  x"13",  x"09", -- 01D0
         x"50",  x"14",  x"09",  x"3a",  x"27",  x"b1",  x"60",  x"47", -- 01D8
         x"2b",  x"3a",  x"26",  x"b1",  x"67",  x"2e",  x"c9",  x"b3", -- 01E0
         x"b4",  x"91",  x"9c",  x"b5",  x"57",  x"88",  x"cd",  x"04", -- 01E8
         x"19",  x"22",  x"c4",  x"9d",  x"21",  x"9d",  x"95",  x"71", -- 01F0
         x"2a",  x"e0",  x"34",  x"07",  x"16",  x"8c",  x"21",  x"ac", -- 01F8
         x"84",  x"49",  x"e3",  x"0e",  x"dc",  x"19",  x"0e",  x"f8", -- 0200
         x"52",  x"c0",  x"32",  x"06",  x"ac",  x"13",  x"1c",  x"21", -- 0208
         x"ba",  x"77",  x"2b",  x"56",  x"1c",  x"60",  x"07",  x"11", -- 0210
         x"28",  x"b1",  x"eb",  x"01",  x"01",  x"73",  x"00",  x"ed", -- 0218
         x"b0",  x"3e",  x"0a",  x"f5",  x"2e",  x"7c",  x"13",  x"7e", -- 0220
         x"00",  x"c6",  x"73",  x"77",  x"23",  x"7e",  x"ce",  x"00", -- 0228
         x"77",  x"50",  x"c3",  x"9c",  x"e1",  x"ad",  x"62",  x"a3", -- 0230
         x"21",  x"44",  x"c8",  x"83",  x"d7",  x"02",  x"d7",  x"00", -- 0238
         x"3e",  x"15",  x"83",  x"4f",  x"37",  x"3e",  x"b2",  x"21", -- 0240
         x"47",  x"52",  x"85",  x"d2",  x"01",  x"c2",  x"7e",  x"02", -- 0248
         x"60",  x"cf",  x"e9",  x"85",  x"83",  x"cf",  x"13",  x"09", -- 0250
         x"7a",  x"c6",  x"09",  x"4f",  x"40",  x"fc",  x"66",  x"d5", -- 0258
         x"48",  x"e5",  x"13",  x"d1",  x"02",  x"14",  x"7a",  x"d6", -- 0260
         x"03",  x"38",  x"e7",  x"70",  x"75",  x"3a",  x"2d",  x"b1", -- 0268
         x"57",  x"cc",  x"56",  x"3a",  x"2c",  x"e4",  x"01",  x"0e", -- 0270
         x"00",  x"7b",  x"b0",  x"32",  x"80",  x"cb",  x"7a",  x"b1", -- 0278
         x"32",  x"c6",  x"80",  x"81",  x"d3",  x"22",  x"81",  x"8e", -- 0280
         x"3a",  x"2f",  x"22",  x"1b",  x"2e",  x"65",  x"1b",  x"28", -- 0288
         x"b4",  x"1b",  x"29",  x"15",  x"31",  x"89",  x"15",  x"30", -- 0290
         x"96",  x"15",  x"2a",  x"15",  x"2b",  x"87",  x"84",  x"8d", -- 0298
         x"21",  x"d0",  x"99",  x"0e",  x"2a",  x"28",  x"ff",  x"4e", -- 02A0
         x"7d",  x"26",  x"28",  x"10",  x"e5",  x"95",  x"0c",  x"66", -- 02A8
         x"8c",  x"03",  x"a8",  x"8d",  x"00",  x"e1",  x"24",  x"7c", -- 02B0
         x"d6",  x"17",  x"38",  x"ef",  x"3e",  x"76",  x"10",  x"1a", -- 02B8
         x"11",  x"3a",  x"e9",  x"69",  x"82",  x"01",  x"b6",  x"20", -- 02C0
         x"12",  x"21",  x"e0",  x"25",  x"59",  x"6d",  x"06",  x"42", -- 02C8
         x"cb",  x"3a",  x"c3",  x"9d",  x"d1",  x"85",  x"e5",  x"b1", -- 02D0
         x"0a",  x"3a",  x"93",  x"02",  x"3d",  x"20",  x"08",  x"21", -- 02D8
         x"f9",  x"84",  x"72",  x"0d",  x"d6",  x"02",  x"89",  x"0e", -- 02E0
         x"00",  x"85",  x"34",  x"0e",  x"ed",  x"93",  x"07",  x"97", -- 02E8
         x"09",  x"64",  x"36",  x"97",  x"03",  x"50",  x"8d",  x"97", -- 02F0
         x"09",  x"92",  x"0e",  x"28",  x"a6",  x"0e",  x"d0",  x"0e", -- 02F8
         x"48",  x"2a",  x"0e",  x"f1",  x"b2",  x"ad",  x"b4",  x"b2", -- 0300
         x"4a",  x"0a",  x"43",  x"dd",  x"68",  x"46",  x"a0",  x"4e", -- 0308
         x"51",  x"ff",  x"fc",  x"81",  x"3c",  x"28",  x"6b",  x"68", -- 0310
         x"61",  x"11",  x"e8",  x"07",  x"a4",  x"21",  x"d0",  x"a9", -- 0318
         x"e5",  x"d5",  x"95",  x"a9",  x"14",  x"c1",  x"aa",  x"92", -- 0320
         x"a2",  x"a6",  x"4e",  x"d0",  x"a6",  x"20",  x"48",  x"db", -- 0328
         x"05",  x"fc",  x"05",  x"42",  x"c7",  x"27",  x"85",  x"26", -- 0330
         x"60",  x"ec",  x"c1",  x"a2",  x"e5",  x"58",  x"c5",  x"ee", -- 0338
         x"4f",  x"09",  x"56",  x"60",  x"09",  x"11",  x"79",  x"1b", -- 0340
         x"47",  x"fa",  x"22",  x"80",  x"89",  x"fa",  x"c1",  x"21", -- 0348
         x"fb",  x"25",  x"80",  x"fb",  x"22",  x"18",  x"8f",  x"7a", -- 0350
         x"16",  x"4f",  x"a7",  x"08",  x"f7",  x"08",  x"10",  x"10", -- 0358
         x"6e",  x"d4",  x"70",  x"f9",  x"8d",  x"e0",  x"c3",  x"4b", -- 0360
         x"43",  x"2d",  x"54",  x"00",  x"41",  x"50",  x"45",  x"20", -- 0368
         x"62",  x"79",  x"20",  x"41",  x"38",  x"46",  x"2e",  x"89", -- 0370
         x"06",  x"42",  x"61",  x"73",  x"69",  x"63",  x"83",  x"e0", -- 0378
         x"0a",  x"4c",  x"61",  x"64",  x"65",  x"c0",  x"02",  x"72", -- 0380
         x"65",  x"73",  x"73",  x"65",  x"3a",  x"c2",  x"15",  x"0a", -- 0388
         x"45",  x"6e",  x"64",  x"24",  x"0d",  x"63",  x"6f",  x"60", -- 0390
         x"70",  x"2d",  x"31",  x"34",  x"2d",  x"31",  x"32",  x"50", -- 0398
         x"38",  x"0d",  x"53",  x"79",  x"73",  x"14",  x"74",  x"65", -- 03A0
         x"6d",  x"32",  x"53",  x"08",  x"74",  x"61",  x"72",  x"74", -- 03A8
         x"a0",  x"33",  x"46",  x"65",  x"68",  x"6c",  x"00",  x"65", -- 03B0
         x"72",  x"21",  x"20",  x"4b",  x"65",  x"69",  x"6e",  x"01", -- 03B8
         x"20",  x"54",  x"61",  x"70",  x"2d",  x"46",  x"69",  x"d3", -- 03C0
         x"0f",  x"df",  x"a4",  x"09",  x"63",  x"e5",  x"06",  x"38", -- 03C8
         x"fb",  x"27",  x"01",  x"6d",  x"89",  x"58",  x"a5",  x"57", -- 03D0
         x"39",  x"4e",  x"0c",  x"d5",  x"e1",  x"21",  x"e4",  x"ff", -- 03D8
         x"39",  x"81",  x"aa",  x"36",  x"ff",  x"53",  x"a4",  x"29", -- 03E0
         x"cf",  x"4a",  x"a8",  x"fc",  x"95",  x"9a",  x"74",  x"fe", -- 03E8
         x"15",  x"fa",  x"9d",  x"c9",  x"fa",  x"c2",  x"fa",  x"29", -- 03F0
         x"80",  x"00",  x"3e",  x"3a",  x"85",  x"5f",  x"3e",  x"b0", -- 03F8
         x"19",  x"8c",  x"57",  x"af",  x"e7",  x"34",  x"0f",  x"c1", -- 0400
         x"db",  x"20",  x"fb",  x"20",  x"fc",  x"1c",  x"cd",  x"05", -- 0408
         x"66",  x"fc",  x"cd",  x"14",  x"d5",  x"95",  x"6c",  x"d1", -- 0410
         x"80",  x"bc",  x"33",  x"86",  x"b8",  x"97",  x"28",  x"b0", -- 0418
         x"d5",  x"c1",  x"4c",  x"cf",  x"a7",  x"f6",  x"4c",  x"7d", -- 0420
         x"d1",  x"e4",  x"54",  x"51",  x"9d",  x"b4",  x"d9",  x"9a", -- 0428
         x"05",  x"fe",  x"95",  x"8a",  x"0a",  x"ba",  x"ae",  x"41", -- 0430
         x"8a",  x"87",  x"a4",  x"dd",  x"69",  x"60",  x"00",  x"c5", -- 0438
         x"af",  x"be",  x"ed",  x"a0",  x"20",  x"fb",  x"c1",  x"a9", -- 0440
         x"09",  x"0a",  x"c1",  x"cc",  x"b8",  x"f3",  x"85",  x"90", -- 0448
         x"fb",  x"fc",  x"55",  x"48",  x"66",  x"fe",  x"30",  x"11", -- 0450
         x"08",  x"65",  x"cb",  x"66",  x"28",  x"10",  x"9b",  x"63", -- 0458
         x"e3",  x"64",  x"f5",  x"c6",  x"ae",  x"f3",  x"98",  x"f2", -- 0460
         x"8b",  x"34",  x"fa",  x"d3",  x"20",  x"0e",  x"da",  x"47", -- 0468
         x"85",  x"d2",  x"22",  x"ff",  x"0d",  x"ed",  x"00",  x"fb", -- 0470
         x"3c",  x"44",  x"49",  x"22",  x"52",  x"3e",  x"41",  x"db", -- 0478
         x"ea",  x"41",  x"db",  x"40",  x"91",  x"01",  x"29",  x"9b", -- 0480
         x"b1",  x"65",  x"26",  x"41",  x"93",  x"61",  x"dc",  x"a8", -- 0488
         x"ec",  x"5a",  x"14",  x"7b",  x"06",  x"dd",  x"96",  x"04", -- 0490
         x"30",  x"1a",  x"9d",  x"a6",  x"4d",  x"44",  x"a4",  x"7c", -- 0498
         x"f1",  x"69",  x"21",  x"c5",  x"00",  x"b1",  x"d1",  x"e1", -- 04A0
         x"df",  x"f5",  x"51",  x"09",  x"38",  x"ea",  x"18",  x"de", -- 04A8
         x"04",  x"4f",  x"21",  x"dd",  x"86",  x"89",  x"d0",  x"d9", -- 04B0
         x"06",  x"fb",  x"f2",  x"4c",  x"7f",  x"06",  x"42",  x"07", -- 04B8
         x"a5",  x"4f",  x"28",  x"34",  x"cf",  x"ba",  x"53",  x"28", -- 04C0
         x"77",  x"80",  x"df",  x"ea",  x"86",  x"44",  x"11",  x"21", -- 04C8
         x"fd",  x"a9",  x"2b",  x"fd",  x"41",  x"24",  x"18",  x"0f", -- 04D0
         x"21",  x"07",  x"87",  x"27",  x"10",  x"06",  x"2a",  x"35", -- 04D8
         x"0d",  x"5e",  x"0e",  x"06",  x"44",  x"4b",  x"17",  x"de", -- 04E0
         x"15",  x"07",  x"47",  x"10",  x"a4",  x"4b",  x"f0",  x"52", -- 04E8
         x"4b",  x"10",  x"39",  x"4b",  x"c9",  x"1c",  x"4a",  x"c3", -- 04F0
         x"2c",  x"c2",  x"8d",  x"d0",  x"92",  x"20",  x"13",  x"e7", -- 04F8
         x"3a",  x"f4",  x"00",  x"2f",  x"52",  x"4f",  x"4d",  x"00", -- 0500
         x"53",  x"2f",  x"42",  x"41",  x"53",  x"49",  x"43",  x"5f", -- 0508
         x"02",  x"43",  x"30",  x"2e",  x"38",  x"37",  x"42",  x"20", -- 0510
         x"9c",  x"e8",  x"fc",  x"8a",  x"4f",  x"6b",  x"05",  x"90", -- 0518
         x"2f",  x"4f",  x"53",  x"88",  x"2c",  x"d4",  x"0a",  x"5f", -- 0520
         x"00",  x"46",  x"96",  x"2c",  x"20",  x"ad",  x"52",  x"f6", -- 0528
         x"1b",  x"89",  x"f7",  x"0a",  x"03",  x"36",  x"f6",  x"01", -- 0530
         x"cd",  x"46",  x"8c",  x"c2",  x"8a",  x"90",  x"36",  x"6f", -- 0538
         x"90",  x"64",  x"2a",  x"22",  x"ad",  x"c5",  x"76",  x"07", -- 0540
         x"86",  x"06",  x"00",  x"b0",  x"86",  x"00",  x"3d",  x"9e", -- 0548
         x"f1",  x"65",  x"7c",  x"cb",  x"de",  x"f6",  x"02",  x"98", -- 0550
         x"8a",  x"4e",  x"13",  x"06",  x"50",  x"f6",  x"1a",  x"16", -- 0558
         x"11",  x"a6",  x"10",  x"d5",  x"ca",  x"c5",  x"31",  x"8f", -- 0560
         x"4b",  x"21",  x"b2",  x"26",  x"ce",  x"14",  x"db",  x"02", -- 0568
         x"01",  x"35",  x"a9",  x"7c",  x"0f",  x"45",  x"07",  x"3e", -- 0570
         x"7c",  x"03",  x"9f",  x"cd",  x"2d",  x"43",  x"86",  x"06", -- 0578
         x"21",  x"96",  x"aa",  x"cf",  x"73",  x"bc",  x"da",  x"61", -- 0580
         x"ba",  x"5a",  x"6f",  x"18",  x"74",  x"a4",  x"25",  x"3e", -- 0588
         x"0c",  x"9b",  x"03",  x"cd",  x"20",  x"fd",  x"20",  x"75", -- 0590
         x"ff",  x"18",  x"10",  x"2f",  x"11",  x"bf",  x"76",  x"81", -- 0598
         x"09",  x"5a",  x"76",  x"18",  x"86",  x"3b",  x"e7",  x"0f", -- 05A0
         x"e7",  x"12",  x"29",  x"8b",  x"40",  x"97",  x"1a",  x"cd", -- 05A8
         x"37",  x"8c",  x"26",  x"f8",  x"85",  x"db",  x"f6",  x"83", -- 05B0
         x"db",  x"fe",  x"df",  x"02",  x"7e",  x"f6",  x"29",  x"45", -- 05B8
         x"9d",  x"e0",  x"07",  x"10",  x"f8",  x"d6",  x"0a",  x"28", -- 05C0
         x"6a",  x"a2",  x"17",  x"c6",  x"ff",  x"b2",  x"be",  x"c2", -- 05C8
         x"0e",  x"0b",  x"ca",  x"c3",  x"88",  x"c2",  x"07",  x"0d", -- 05D0
         x"ca",  x"19",  x"89",  x"c5",  x"07",  x"1b",  x"28",  x"42", -- 05D8
         x"89",  x"06",  x"1f",  x"ca",  x"d1",  x"04",  x"0e",  x"20", -- 05E0
         x"ca",  x"15",  x"82",  x"07",  x"42",  x"ca",  x"f3",  x"40", -- 05E8
         x"26",  x"44",  x"ca",  x"1e",  x"8a",  x"b1",  x"07",  x"52", -- 05F0
         x"ca",  x"6b",  x"20",  x"07",  x"62",  x"28",  x"72",  x"b4", -- 05F8
         x"06",  x"64",  x"ca",  x"16",  x"72",  x"16",  x"14",  x"c3", -- 0600
         x"73",  x"8a",  x"d4",  x"20",  x"cd",  x"d8",  x"8d",  x"c3", -- 0608
         x"84",  x"fc",  x"13",  x"69",  x"e7",  x"cf",  x"30",  x"0f", -- 0610
         x"06",  x"6e",  x"14",  x"96",  x"f6",  x"da",  x"0f",  x"34", -- 0618
         x"54",  x"f6",  x"15",  x"a1",  x"cc",  x"63",  x"fd",  x"ab", -- 0620
         x"0f",  x"f7",  x"0f",  x"ec",  x"0a",  x"1d",  x"29",  x"30", -- 0628
         x"09",  x"c2",  x"70",  x"94",  x"bd",  x"1f",  x"08",  x"f7", -- 0630
         x"ed",  x"e3",  x"7e",  x"06",  x"20",  x"f5",  x"95",  x"35", -- 0638
         x"f7",  x"0d",  x"40",  x"bd",  x"fc",  x"4c",  x"85",  x"83", -- 0640
         x"34",  x"1f",  x"21",  x"10",  x"75",  x"8b",  x"e5",  x"96", -- 0648
         x"d9",  x"48",  x"0e",  x"e6",  x"e2",  x"d2",  x"f0",  x"41", -- 0650
         x"fd",  x"55",  x"01",  x"e5",  x"e3",  x"e1",  x"28",  x"d6", -- 0658
         x"98",  x"49",  x"ad",  x"d6",  x"df",  x"f5",  x"13",  x"85", -- 0660
         x"8b",  x"52",  x"0c",  x"fa",  x"ca",  x"ed",  x"d2",  x"b6", -- 0668
         x"df",  x"f3",  x"da",  x"fa",  x"66",  x"07",  x"77",  x"fb", -- 0670
         x"f7",  x"c3",  x"dd",  x"8e",  x"fc",  x"07",  x"a9",  x"c4", -- 0678
         x"a7",  x"0d",  x"f9",  x"05",  x"4a",  x"0b",  x"fa",  x"37", -- 0680
         x"db",  x"f1",  x"0b",  x"25",  x"46",  x"fa",  x"3a",  x"a4", -- 0688
         x"0e",  x"e3",  x"56",  x"d0",  x"4a",  x"b5",  x"ca",  x"11", -- 0690
         x"a9",  x"76",  x"7e",  x"f4",  x"22",  x"34",  x"21",  x"87", -- 0698
         x"50",  x"98",  x"a7",  x"24",  x"11",  x"78",  x"2b",  x"f9", -- 06A0
         x"51",  x"e8",  x"49",  x"13",  x"39",  x"f0",  x"a3",  x"af", -- 06A8
         x"82",  x"cc",  x"aa",  x"c4",  x"9f",  x"b5",  x"14",  x"c9", -- 06B0
         x"d5",  x"ca",  x"aa",  x"97",  x"33",  x"a4",  x"10",  x"30", -- 06B8
         x"60",  x"74",  x"69",  x"5d",  x"cb",  x"7b",  x"20",  x"13", -- 06C0
         x"ab",  x"0c",  x"d4",  x"d0",  x"d6",  x"2f",  x"20",  x"03", -- 06C8
         x"e9",  x"87",  x"05",  x"81",  x"cf",  x"1d",  x"18",  x"ea", -- 06D0
         x"da",  x"8b",  x"4e",  x"64",  x"19",  x"34",  x"88",  x"21", -- 06D8
         x"32",  x"5e",  x"18",  x"66",  x"5d",  x"b7",  x"31",  x"ed", -- 06E0
         x"5b",  x"9a",  x"67",  x"3a",  x"06",  x"93",  x"3a",  x"bf", -- 06E8
         x"e2",  x"9a",  x"30",  x"52",  x"6e",  x"f3",  x"27",  x"26", -- 06F0
         x"20",  x"93",  x"ea",  x"10",  x"55",  x"46",  x"f0",  x"1f", -- 06F8
         x"34",  x"20",  x"e5",  x"ed",  x"20",  x"34",  x"a7",  x"ec", -- 0700
         x"db",  x"ef",  x"96",  x"80",  x"ee",  x"80",  x"d6",  x"90", -- 0708
         x"38",  x"e2",  x"9d",  x"c1",  x"0b",  x"18",  x"b9",  x"d6", -- 0710
         x"2d",  x"bd",  x"0a",  x"18",  x"11",  x"e9",  x"28",  x"eb", -- 0718
         x"86",  x"ca",  x"e6",  x"35",  x"ae",  x"00",  x"c3",  x"0d", -- 0720
         x"88",  x"46",  x"53",  x"20",  x"74",  x"67",  x"96",  x"6f", -- 0728
         x"3a",  x"75",  x"6e",  x"9c",  x"6d",  x"74",  x"8e",  x"52", -- 0730
         x"0d",  x"b4",  x"aa",  x"b5",  x"e9",  x"d6",  x"a1",  x"16", -- 0738
         x"72",  x"2e",  x"6f",  x"6c",  x"de",  x"87",  x"53",  x"44", -- 0740
         x"43",  x"ef",  x"43",  x"64",  x"20",  x"6b",  x"11",  x"a3", -- 0748
         x"29",  x"20",  x"6e",  x"e9",  x"62",  x"68",  x"74",  x"81", -- 0750
         x"38",  x"6f",  x"65",  x"66",  x"66",  x"6e",  x"9e",  x"38", -- 0758
         x"20",  x"77",  x"31",  x"d1",  x"ca",  x"6e",  x"d9",  x"60", -- 0760
         x"2a",  x"20",  x"43",  x"75",  x"15",  x"72",  x"73",  x"6f", -- 0768
         x"99",  x"7d",  x"ed",  x"78",  x"10",  x"38",  x"4e",  x"61", -- 0770
         x"76",  x"06",  x"69",  x"67",  x"61",  x"74",  x"69",  x"36", -- 0778
         x"0a",  x"dd",  x"1a",  x"45",  x"3a",  x"83",  x"59",  x"41", -- 0780
         x"75",  x"73",  x"77",  x"61",  x"64",  x"a0",  x"10",  x"53", -- 0788
         x"70",  x"61",  x"63",  x"ab",  x"89",  x"1a",  x"49",  x"6e", -- 0790
         x"66",  x"31",  x"6d",  x"5a",  x"25",  x"41",  x"64",  x"42", -- 0798
         x"14",  x"6b",  x"73",  x"ac",  x"19",  x"56",  x"2f",  x"7a", -- 07A0
         x"65",  x"ac",  x"6b",  x"6f",  x"73",  x"20",  x"3b",  x"68", -- 07A8
         x"6f",  x"07",  x"44",  x"c3",  x"95",  x"17",  x"6f",  x"76", -- 07B0
         x"17",  x"6c",  x"61",  x"f8",  x"bb",  x"55",  x"25",  x"42", -- 07B8
         x"3a",  x"fa",  x"73",  x"2d",  x"50",  x"aa",  x"00",  x"67", -- 07C0
         x"72",  x"61",  x"6d",  x"17",  x"6d",  x"20",  x"73",  x"9a", -- 07C8
         x"95",  x"1b",  x"84",  x"b5",  x"b2",  x"09",  x"fb",  x"1f", -- 07D0
         x"26",  x"ed",  x"8f",  x"00",  x"43",  x"44",  x"15",  x"03", -- 07D8
         x"15",  x"20",  x"55",  x"70",  x"0d",  x"f7",  x"bc",  x"3c", -- 07E0
         x"30",  x"d6",  x"37",  x"56",  x"fa",  x"0a",  x"30",  x"30", -- 07E8
         x"31",  x"20",  x"11",  x"c5",  x"1e",  x"db",  x"00",  x"b7", -- 07F0
         x"1b",  x"8e",  x"02",  x"98",  x"a0",  x"7e",  x"d3",  x"00", -- 07F8
         x"c9",  x"33",  x"db",  x"01",  x"af",  x"00",  x"02",  x"d3", -- 0800
         x"01",  x"6f",  x"c9",  x"c1",  x"e1",  x"e5",  x"66",  x"c5", -- 0808
         x"bb",  x"c8",  x"25",  x"23",  x"e5",  x"ca",  x"10",  x"e1", -- 0810
         x"18",  x"f2",  x"c9",  x"50",  x"fd",  x"24",  x"fd",  x"39", -- 0818
         x"fd",  x"66",  x"56",  x"04",  x"7e",  x"00",  x"af",  x"c0", -- 0820
         x"30",  x"0a",  x"7a",  x"c6",  x"30",  x"95",  x"1c",  x"c9", -- 0828
         x"a6",  x"09",  x"37",  x"09",  x"91",  x"47",  x"07",  x"45", -- 0830
         x"00",  x"e6",  x"0f",  x"39",  x"11",  x"d3",  x"11",  x"27", -- 0838
         x"10",  x"0c",  x"9c",  x"42",  x"66",  x"01",  x"7f",  x"2e", -- 0840
         x"9d",  x"21",  x"aa",  x"4f",  x"10",  x"36",  x"0e",  x"3f", -- 0848
         x"25",  x"18",  x"00",  x"56",  x"7a",  x"82",  x"2b",  x"05", -- 0850
         x"07",  x"d5",  x"36",  x"6a",  x"0e",  x"2c",  x"7c",  x"b2", -- 0858
         x"06",  x"f1",  x"00",  x"ec",  x"36",  x"20",  x"5d",  x"54", -- 0860
         x"13",  x"01",  x"3f",  x"bf",  x"03",  x"8a",  x"d1",  x"0c", -- 0868
         x"e8",  x"32",  x"0c",  x"b4",  x"6e",  x"32",  x"24",  x"c9", -- 0870
         x"f2",  x"c4",  x"ed",  x"67",  x"4b",  x"0c",  x"06",  x"00", -- 0878
         x"d5",  x"9a",  x"c2",  x"a9",  x"09",  x"c6",  x"5f",  x"11", -- 0880
         x"2c",  x"aa",  x"a6",  x"5e",  x"04",  x"ca",  x"67",  x"d5", -- 0888
         x"01",  x"28",  x"4a",  x"a8",  x"1e",  x"d3",  x"be",  x"00", -- 0890
         x"ee",  x"d9",  x"08",  x"50",  x"2d",  x"20",  x"9a",  x"2d", -- 0898
         x"3b",  x"3c",  x"2e",  x"ec",  x"19",  x"c3",  x"88",  x"84", -- 08A0
         x"66",  x"04",  x"84",  x"ca",  x"05",  x"da",  x"d2",  x"4a", -- 08A8
         x"03",  x"b4",  x"d8",  x"d6",  x"09",  x"29",  x"28",  x"21", -- 08B0
         x"d5",  x"f1",  x"9d",  x"6b",  x"20",  x"f4",  x"b4",  x"2b", -- 08B8
         x"34",  x"e0",  x"f3",  x"04",  x"4e",  x"6b",  x"62",  x"2c", -- 08C0
         x"44",  x"19",  x"10",  x"30",  x"18",  x"d3",  x"8d",  x"15", -- 08C8
         x"b5",  x"a8",  x"28",  x"19",  x"b9",  x"3a",  x"12",  x"13", -- 08D0
         x"05",  x"18",  x"b2",  x"3e",  x"17",  x"fd",  x"02",  x"3d", -- 08D8
         x"fd",  x"96",  x"00",  x"30",  x"05",  x"41",  x"80",  x"43", -- 08E0
         x"33",  x"a0",  x"84",  x"01",  x"7b",  x"12",  x"f8",  x"7f", -- 08E8
         x"c1",  x"b1",  x"3d",  x"04",  x"e8",  x"62",  x"4f",  x"47", -- 08F0
         x"1b",  x"79",  x"47",  x"88",  x"9e",  x"07",  x"78",  x"c8", -- 08F8
         x"9e",  x"77",  x"eb",  x"db",  x"9c",  x"06",  x"6c",  x"37", -- 0900
         x"06",  x"06",  x"a4",  x"06",  x"cb",  x"05",  x"3e",  x"03", -- 0908
         x"04",  x"3a",  x"1e",  x"10",  x"82",  x"2c",  x"34",  x"ff", -- 0910
         x"a2",  x"05",  x"04",  x"38",  x"cf",  x"c2",  x"57",  x"26", -- 0918
         x"4e",  x"06",  x"28",  x"e0",  x"20",  x"23",  x"10",  x"fb", -- 0920
         x"c9",  x"01",  x"28",  x"07",  x"00",  x"0e",  x"21",  x"d0", -- 0928
         x"62",  x"8d",  x"e7",  x"c3",  x"ce",  x"07",  x"3e",  x"05", -- 0930
         x"9c",  x"f2",  x"06",  x"f0",  x"c9",  x"aa",  x"ca",  x"cd", -- 0938
         x"0a",  x"31",  x"00",  x"0d",  x"89",  x"d8",  x"0d",  x"0a", -- 0940
         x"c1",  x"d1",  x"ed",  x"03",  x"53",  x"d7",  x"03",  x"21", -- 0948
         x"bd",  x"c0",  x"2d",  x"0c",  x"03",  x"01",  x"67",  x"00", -- 0950
         x"2d",  x"eb",  x"f9",  x"00",  x"af",  x"32",  x"ab",  x"03", -- 0958
         x"32",  x"00",  x"04",  x"2a",  x"50",  x"36",  x"41",  x"ff", -- 0960
         x"22",  x"b0",  x"03",  x"03",  x"19",  x"22",  x"56",  x"03", -- 0968
         x"3e",  x"14",  x"00",  x"fc",  x"03",  x"cd",  x"4f",  x"c6", -- 0970
         x"23",  x"eb",  x"cd",  x"00",  x"93",  x"c4",  x"cd",  x"69", -- 0978
         x"c6",  x"c3",  x"54",  x"c8",  x"42",  x"c9",  x"42",  x"3a", -- 0980
         x"21",  x"c0",  x"01",  x"aa",  x"2c",  x"1f",  x"12",  x"42", -- 0988
         x"d7",  x"41",  x"5e",  x"41",  x"21",  x"49",  x"31",  x"67", -- 0990
         x"75",  x"24",  x"0d",  x"60",  x"47",  x"3e",  x"ff",  x"d3", -- 0998
         x"04",  x"db",  x"52",  x"05",  x"c6",  x"0c",  x"db",  x"04", -- 09A0
         x"6f",  x"0c",  x"3c",  x"d3",  x"4a",  x"07",  x"98",  x"75", -- 09A8
         x"07",  x"27",  x"15",  x"c8",  x"40",  x"d3",  x"06",  x"c3", -- 09B0
         x"6d",  x"8e",  x"93",  x"0b",  x"09",  x"96",  x"13",  x"50", -- 09B8
         x"20",  x"04",  x"c9",  x"16",  x"5a",  x"44",  x"00",  x"9a", -- 09C0
         x"00",  x"15",  x"7a",  x"19",  x"f0",  x"20",  x"ea",  x"68", -- 09C8
         x"ae",  x"54",  x"7e",  x"ce",  x"5b",  x"05",  x"be",  x"af", -- 09D0
         x"16",  x"09",  x"c0",  x"94",  x"13",  x"e5",  x"b2",  x"03", -- 09D8
         x"3e",  x"77",  x"90",  x"cc",  x"bb",  x"8e",  x"a3",  x"9b", -- 09E0
         x"c3",  x"57",  x"95",  x"da",  x"97",  x"8f",  x"ce",  x"05", -- 09E8
         x"8e",  x"0d",  x"f9",  x"07",  x"13",  x"9b",  x"8e",  x"33", -- 09F0
         x"f5",  x"f5",  x"2e",  x"05",  x"fb",  x"43",  x"06",  x"dd", -- 09F8
         x"56",  x"07",  x"c8",  x"30",  x"08",  x"f1",  x"06",  x"18", -- 0A00
         x"00",  x"cb",  x"3b",  x"cb",  x"1a",  x"cb",  x"1d",  x"cb", -- 0A08
         x"1c",  x"c5",  x"f5",  x"e5",  x"09",  x"a1",  x"1f",  x"10", -- 0A10
         x"e4",  x"1f",  x"08",  x"7d",  x"1f",  x"4a",  x"1e",  x"08", -- 0A18
         x"26",  x"50",  x"01",  x"73",  x"d6",  x"40",  x"20",  x"16", -- 0A20
         x"02",  x"26",  x"95",  x"08",  x"48",  x"a4",  x"08",  x"87", -- 0A28
         x"a7",  x"19",  x"16",  x"0a",  x"b2",  x"58",  x"eb",  x"0d", -- 0A30
         x"d1",  x"cb",  x"7d",  x"c4",  x"6c",  x"ce",  x"14",  x"f2", -- 0A38
         x"bb",  x"1a",  x"9c",  x"34",  x"08",  x"cd",  x"28",  x"87", -- 0A40
         x"8e",  x"a8",  x"11",  x"e1",  x"46",  x"c9",  x"f5",  x"01", -- 0A48
         x"f5",  x"3b",  x"cd",  x"7a",  x"8e",  x"26",  x"64",  x"b5", -- 0A50
         x"1a",  x"a8",  x"17",  x"25",  x"73",  x"dd",  x"f6",  x"b4", -- 0A58
         x"ab",  x"26",  x"96",  x"0b",  x"cf",  x"d0",  x"df",  x"08", -- 0A60
         x"a0",  x"f5",  x"4e",  x"40",  x"f5",  x"01",  x"2d",  x"c2", -- 0A68
         x"24",  x"91",  x"2a",  x"4d",  x"af",  x"63",  x"1e",  x"aa", -- 0A70
         x"01",  x"1e",  x"44",  x"48",  x"94",  x"1e",  x"ac",  x"90", -- 0A78
         x"15",  x"39",  x"cc",  x"f3",  x"00",  x"68",  x"f1",  x"cc", -- 0A80
         x"19",  x"bd",  x"c5",  x"81",  x"8e",  x"7d",  x"d1",  x"b8", -- 0A88
         x"cf",  x"77",  x"04",  x"78",  x"a3",  x"f4",  x"25",  x"eb", -- 0A90
         x"d5",  x"3b",  x"68",  x"d1",  x"ff",  x"23",  x"14",  x"23", -- 0A98
         x"7e",  x"3d",  x"4b",  x"d5",  x"37",  x"fd",  x"e1",  x"d0", -- 0AA0
         x"14",  x"03",  x"d6",  x"aa",  x"0a",  x"01",  x"03",  x"10", -- 0AA8
         x"27",  x"78",  x"b1",  x"28",  x"28",  x"32",  x"95",  x"79", -- 0AB0
         x"40",  x"2a",  x"79",  x"e9",  x"7a",  x"5a",  x"45",  x"c1", -- 0AB8
         x"ca",  x"0a",  x"58",  x"50",  x"b0",  x"63",  x"09",  x"0b", -- 0AC0
         x"18",  x"d4",  x"2b",  x"52",  x"ca",  x"3e",  x"af",  x"28", -- 0AC8
         x"a4",  x"11",  x"7a",  x"2a",  x"2a",  x"b7",  x"4f",  x"42", -- 0AD0
         x"47",  x"81",  x"81",  x"88",  x"d1",  x"77",  x"28",  x"04", -- 0AD8
         x"ec",  x"92",  x"18",  x"02",  x"29",  x"3e",  x"04",  x"b2", -- 0AE0
         x"9c",  x"c3",  x"26",  x"60",  x"e7",  x"22",  x"e9",  x"88", -- 0AE8
         x"dd",  x"38",  x"08",  x"a1",  x"86",  x"05",  x"02",  x"16", -- 0AF0
         x"e9",  x"18",  x"06",  x"09",  x"07",  x"01",  x"16",  x"41", -- 0AF8
         x"41",  x"9f",  x"26",  x"c5",  x"50",  x"a1",  x"31",  x"d5", -- 0B00
         x"50",  x"9d",  x"52",  x"d6",  x"29",  x"1a",  x"25",  x"27", -- 0B08
         x"02",  x"a2",  x"59",  x"50",  x"03",  x"9c",  x"27",  x"4a", -- 0B10
         x"04",  x"b0",  x"c1",  x"ff",  x"32",  x"1f",  x"b2",  x"42", -- 0B18
         x"8f",  x"3e",  x"52",  x"02",  x"1a",  x"7f",  x"8b",  x"de", -- 0B20
         x"10",  x"ae",  x"1a",  x"9b",  x"70",  x"9a",  x"64",  x"2e", -- 0B28
         x"df",  x"f9",  x"8b",  x"ab",  x"23",  x"3b",  x"21",  x"28", -- 0B30
         x"06",  x"cb",  x"5e",  x"20",  x"16",  x"f5",  x"94",  x"7b", -- 0B38
         x"eb",  x"0c",  x"cb",  x"06",  x"26",  x"03",  x"07",  x"16", -- 0B40
         x"d4",  x"03",  x"08",  x"03",  x"09",  x"15",  x"16",  x"10", -- 0B48
         x"ee",  x"4c",  x"7b",  x"e1",  x"9e",  x"b9",  x"af",  x"02", -- 0B50
         x"66",  x"09",  x"e5",  x"cc",  x"c0",  x"66",  x"07",  x"d1", -- 0B58
         x"6f",  x"51",  x"20",  x"6f",  x"20",  x"74",  x"11",  x"40", -- 0B60
         x"9c",  x"90",  x"97",  x"c0",  x"7d",  x"3c",  x"20",  x"05", -- 0B68
         x"1b",  x"7a",  x"66",  x"b3",  x"97",  x"7d",  x"0c",  x"d6", -- 0B70
         x"fe",  x"20",  x"5e",  x"78",  x"dd",  x"96",  x"28",  x"0a", -- 0B78
         x"67",  x"05",  x"9e",  x"0b",  x"31",  x"6f",  x"7c",  x"0a", -- 0B80
         x"0c",  x"67",  x"7d",  x"bf",  x"09",  x"0d",  x"f9",  x"62", -- 0B88
         x"fd",  x"97",  x"fe",  x"c0",  x"8b",  x"0b",  x"dd",  x"0d", -- 0B90
         x"b6",  x"0a",  x"28",  x"10",  x"4d",  x"0a",  x"94",  x"4d", -- 0B98
         x"0b",  x"e5",  x"3b",  x"e1",  x"19",  x"2b",  x"7c",  x"b5", -- 0BA0
         x"98",  x"eb",  x"0f",  x"04",  x"a4",  x"43",  x"5e",  x"0c", -- 0BA8
         x"a4",  x"42",  x"0d",  x"e5",  x"51",  x"d9",  x"c5",  x"d8", -- 0BB0
         x"23",  x"6e",  x"52",  x"f1",  x"b2",  x"e2",  x"a8",  x"26", -- 0BB8
         x"df",  x"28",  x"d9",  x"34",  x"2d",  x"ff",  x"60",  x"c8", -- 0BC0
         x"4e",  x"3d",  x"08",  x"c7",  x"3d",  x"09",  x"43",  x"4a", -- 0BC8
         x"a9",  x"03",  x"b0",  x"28",  x"07",  x"68",  x"7d",  x"06", -- 0BD0
         x"3f",  x"de",  x"c6",  x"25",  x"99",  x"24",  x"d3",  x"81", -- 0BD8
         x"82",  x"e5",  x"29",  x"a0",  x"5b",  x"1f",  x"05",  x"fc", -- 0BE0
         x"05",  x"cb",  x"28",  x"77",  x"fd",  x"1e",  x"60",  x"4e", -- 0BE8
         x"3b",  x"46",  x"09",  x"51",  x"58",  x"0b",  x"0f",  x"7b", -- 0BF0
         x"b2",  x"28",  x"2e",  x"4e",  x"24",  x"1c",  x"66",  x"ff", -- 0BF8
         x"7e",  x"d2",  x"60",  x"cb",  x"03",  x"a8",  x"d7",  x"0c", -- 0C00
         x"5f",  x"17",  x"9f",  x"57",  x"84",  x"29",  x"0e",  x"fc", -- 0C08
         x"66",  x"0e",  x"fd",  x"67",  x"0e",  x"6f",  x"00",  x"7b", -- 0C10
         x"94",  x"5f",  x"7a",  x"9d",  x"57",  x"6b",  x"7a",  x"08", -- 0C18
         x"67",  x"b3",  x"28",  x"cb",  x"c0",  x"89",  x"07",  x"21", -- 0C20
         x"ef",  x"ff",  x"39",  x"f9",  x"8a",  x"45",  x"20",  x"b2", -- 0C28
         x"aa",  x"bf",  x"02",  x"9f",  x"6a",  x"de",  x"14",  x"69", -- 0C30
         x"6c",  x"04",  x"07",  x"04",  x"38",  x"21",  x"b4",  x"95", -- 0C38
         x"00",  x"66",  x"06",  x"fd",  x"6e",  x"07",  x"fd",  x"46", -- 0C40
         x"08",  x"14",  x"fd",  x"4e",  x"09",  x"24",  x"94",  x"a5", -- 0C48
         x"23",  x"9d",  x"28",  x"22",  x"98",  x"21",  x"99",  x"38", -- 0C50
         x"1c",  x"09",  x"21",  x"01",  x"99",  x"60",  x"47",  x"c3", -- 0C58
         x"3d",  x"95",  x"1a",  x"67",  x"00",  x"d6",  x"01",  x"da", -- 0C60
         x"37",  x"95",  x"3e",  x"03",  x"94",  x"a1",  x"05",  x"7c", -- 0C68
         x"c6",  x"ff",  x"61",  x"b2",  x"25",  x"94",  x"d7",  x"9e", -- 0C70
         x"b4",  x"19",  x"ee",  x"14",  x"c5",  x"21",  x"10",  x"8c", -- 0C78
         x"a5",  x"01",  x"04",  x"43",  x"dd",  x"c1",  x"f7",  x"07", -- 0C80
         x"ff",  x"f8",  x"41",  x"21",  x"22",  x"93",  x"19",  x"80", -- 0C88
         x"00",  x"d1",  x"e9",  x"c3",  x"2b",  x"93",  x"c3",  x"40", -- 0C90
         x"0e",  x"94",  x"c3",  x"b8",  x"94",  x"fc",  x"4d",  x"cb", -- 0C98
         x"3c",  x"e4",  x"80",  x"09",  x"4d",  x"7c",  x"e6",  x"01", -- 0CA0
         x"47",  x"1b",  x"7c",  x"cb",  x"3f",  x"3f",  x"f7",  x"bc", -- 0CA8
         x"13",  x"f8",  x"00",  x"03",  x"52",  x"f9",  x"03",  x"fa", -- 0CB0
         x"80",  x"8f",  x"fb",  x"dd",  x"67",  x"86",  x"11",  x"77", -- 0CB8
         x"f3",  x"08",  x"89",  x"84",  x"8e",  x"f8",  x"b6",  x"08", -- 0CC0
         x"f4",  x"08",  x"fd",  x"08",  x"f9",  x"e8",  x"08",  x"a5", -- 0CC8
         x"5b",  x"fe",  x"08",  x"fa",  x"08",  x"32",  x"f6",  x"79", -- 0CD0
         x"d4",  x"d0",  x"da",  x"3d",  x"28",  x"48",  x"2c",  x"f7", -- 0CD8
         x"b5",  x"d9",  x"1a",  x"f2",  x"63",  x"98",  x"4f",  x"ca", -- 0CE0
         x"bf",  x"b4",  x"06",  x"94",  x"36",  x"66",  x"f4",  x"a6", -- 0CE8
         x"46",  x"46",  x"91",  x"bb",  x"2b",  x"0a",  x"e9",  x"d6", -- 0CF0
         x"f9",  x"8c",  x"67",  x"ca",  x"1e",  x"75",  x"85",  x"a9", -- 0CF8
         x"8c",  x"2b",  x"4d",  x"44",  x"c5",  x"e6",  x"34",  x"b1", -- 0D00
         x"a0",  x"ca",  x"d3",  x"a1",  x"c1",  x"34",  x"e5",  x"69", -- 0D08
         x"34",  x"fd",  x"e5",  x"17",  x"35",  x"48",  x"dc",  x"c2", -- 0D10
         x"c2",  x"34",  x"eb",  x"5e",  x"23",  x"56",  x"98",  x"b6", -- 0D18
         x"2b",  x"6e",  x"28",  x"67",  x"7b",  x"94",  x"31",  x"d9", -- 0D20
         x"a0",  x"90",  x"28",  x"57",  x"7d",  x"8c",  x"28",  x"bc", -- 0D28
         x"f0",  x"88",  x"06",  x"67",  x"1c",  x"20",  x"07",  x"14", -- 0D30
         x"88",  x"00",  x"2c",  x"20",  x"01",  x"24",  x"03",  x"a6", -- 0D38
         x"57",  x"01",  x"55",  x"c5",  x"fe",  x"02",  x"03",  x"7d", -- 0D40
         x"36",  x"49",  x"ec",  x"47",  x"7c",  x"7e",  x"23",  x"2a", -- 0D48
         x"66",  x"6f",  x"dc",  x"5a",  x"46",  x"b3",  x"f9",  x"9d", -- 0D50
         x"62",  x"80",  x"10",  x"18",  x"fa",  x"18",  x"04",  x"82", -- 0D58
         x"92",  x"0f",  x"67",  x"8b",  x"d5",  x"69",  x"b9",  x"62", -- 0D60
         x"29",  x"eb",  x"83",  x"8e",  x"c8",  x"16",  x"6e",  x"84", -- 0D68
         x"6c",  x"46",  x"81",  x"cd",  x"4e",  x"07",  x"90",  x"b9", -- 0D70
         x"8e",  x"17",  x"39",  x"cb",  x"18",  x"8e",  x"27",  x"3d", -- 0D78
         x"20",  x"19",  x"8a",  x"96",  x"84",  x"51",  x"94",  x"4a", -- 0D80
         x"8d",  x"92",  x"29",  x"88",  x"45",  x"90",  x"89",  x"43", -- 0D88
         x"8e",  x"12",  x"da",  x"16",  x"8b",  x"28",  x"d5",  x"6c", -- 0D90
         x"d6",  x"24",  x"d5",  x"0c",  x"80",  x"ac",  x"8b",  x"26", -- 0D98
         x"77",  x"2a",  x"cb",  x"bd",  x"79",  x"10",  x"7a",  x"41", -- 0DA0
         x"07",  x"8a",  x"7a",  x"04",  x"08",  x"0f",  x"7a",  x"20", -- 0DA8
         x"11",  x"79",  x"ce",  x"13",  x"46",  x"23",  x"d4",  x"10", -- 0DB0
         x"4e",  x"6a",  x"60",  x"79",  x"c1",  x"fa",  x"57",  x"bc", -- 0DB8
         x"e7",  x"a7",  x"d5",  x"1a",  x"fb",  x"c9",  x"f5",  x"90", -- 0DC0
         x"a5",  x"c6",  x"fe",  x"d4",  x"60",  x"04",  x"84",  x"8a", -- 0DC8
         x"ce",  x"e2",  x"35",  x"05",  x"25",  x"88",  x"a9",  x"07", -- 0DD0
         x"06",  x"8c",  x"2d",  x"07",  x"07",  x"69",  x"af",  x"b6", -- 0DD8
         x"f7",  x"b2",  x"93",  x"23",  x"af",  x"7d",  x"2c",  x"cb", -- 0DE0
         x"93",  x"18",  x"33",  x"67",  x"78",  x"03",  x"47",  x"79", -- 0DE8
         x"03",  x"52",  x"4f",  x"3e",  x"95",  x"91",  x"3a",  x"9c", -- 0DF0
         x"08",  x"bf",  x"07",  x"aa",  x"5b",  x"f2",  x"f5",  x"4e", -- 0DF8
         x"d3",  x"86",  x"4e",  x"aa",  x"aa",  x"0d",  x"67",  x"d5", -- 0E00
         x"b5",  x"33",  x"b9",  x"ca",  x"a4",  x"d8",  x"ac",  x"0a", -- 0E08
         x"52",  x"a8",  x"f1",  x"00",  x"32",  x"dd",  x"72",  x"5f", -- 0E10
         x"73",  x"fe",  x"dc",  x"94",  x"75",  x"fc",  x"3f",  x"e1", -- 0E18
         x"11",  x"eb",  x"2c",  x"19",  x"56",  x"b0",  x"30",  x"b6", -- 0E20
         x"a0",  x"ff",  x"28",  x"82",  x"6f",  x"fd",  x"0b",  x"8b", -- 0E28
         x"67",  x"fb",  x"05",  x"5f",  x"41",  x"bb",  x"88",  x"57", -- 0E30
         x"1c",  x"b8",  x"0c",  x"2a",  x"b7",  x"28",  x"cd",  x"28", -- 0E38
         x"84",  x"c1",  x"7e",  x"d6",  x"03",  x"20",  x"1f",  x"60", -- 0E40
         x"c2",  x"14",  x"58",  x"6f",  x"c0",  x"14",  x"00",  x"67", -- 0E48
         x"c7",  x"74",  x"16",  x"3e",  x"f4",  x"80",  x"23",  x"cb", -- 0E50
         x"04",  x"12",  x"cb",  x"11",  x"cb",  x"10",  x"83",  x"d6", -- 0E58
         x"a6",  x"1e",  x"1a",  x"1e",  x"c9",  x"8f",  x"6e",  x"6c", -- 0E60
         x"f3",  x"75",  x"c5",  x"73",  x"36",  x"fe",  x"00",  x"be", -- 0E68
         x"ca",  x"ee",  x"61",  x"b6",  x"fc",  x"6f",  x"7a",  x"ec", -- 0E70
         x"04",  x"d3",  x"79",  x"c6",  x"04",  x"fe",  x"5f",  x"78", -- 0E78
         x"04",  x"ff",  x"8f",  x"6c",  x"91",  x"6e",  x"e3",  x"2a", -- 0E80
         x"fa",  x"e2",  x"d7",  x"af",  x"dc",  x"d3",  x"77",  x"c5", -- 0E88
         x"bb",  x"d9",  x"a7",  x"c8",  x"2d",  x"fa",  x"fd",  x"c8", -- 0E90
         x"dd",  x"fb",  x"05",  x"bf",  x"c8",  x"05",  x"6f",  x"c8", -- 0E98
         x"b5",  x"66",  x"fa",  x"72",  x"12",  x"16",  x"c9",  x"84", -- 0EA0
         x"4a",  x"0c",  x"c8",  x"0f",  x"05",  x"1a",  x"c3",  x"c9", -- 0EA8
         x"fb",  x"96",  x"21",  x"bd",  x"e4",  x"11",  x"06",  x"a1", -- 0EB0
         x"e1",  x"49",  x"e5",  x"49",  x"9f",  x"a9",  x"26",  x"92", -- 0EB8
         x"24",  x"9b",  x"4a",  x"22",  x"9c",  x"20",  x"1d",  x"9d", -- 0EC0
         x"38",  x"05",  x"98",  x"0c",  x"c3",  x"64",  x"97",  x"0a", -- 0EC8
         x"f8",  x"c6",  x"50",  x"0e",  x"f1",  x"30",  x"f9",  x"aa", -- 0ED0
         x"55",  x"57",  x"16",  x"06",  x"9b",  x"02",  x"fb",  x"c7", -- 0ED8
         x"02",  x"fa",  x"20",  x"15",  x"3f",  x"60",  x"ea",  x"0e", -- 0EE0
         x"a6",  x"f5",  x"e7",  x"46",  x"f5",  x"60",  x"d1",  x"21", -- 0EE8
         x"08",  x"00",  x"6b",  x"09",  x"11",  x"eb",  x"12",  x"9d", -- 0EF0
         x"11",  x"0c",  x"e1",  x"11",  x"dd",  x"42",  x"d4",  x"ff", -- 0EF8
         x"8b",  x"3e",  x"31",  x"28",  x"17",  x"f9",  x"d9",  x"0a", -- 0F00
         x"66",  x"a6",  x"ed",  x"06",  x"fa",  x"06",  x"fb",  x"91", -- 0F08
         x"80",  x"42",  x"95",  x"8e",  x"fe",  x"cd",  x"61",  x"18", -- 0F10
         x"08",  x"eb",  x"4e",  x"21",  x"a5",  x"a5",  x"56",  x"ee", -- 0F18
         x"80",  x"71",  x"23",  x"70",  x"23",  x"1d",  x"73",  x"23", -- 0F20
         x"72",  x"a6",  x"c6",  x"c2",  x"cf",  x"f0",  x"a2",  x"cf", -- 0F28
         x"c6",  x"81",  x"32",  x"bb",  x"64",  x"30",  x"a6",  x"39", -- 0F30
         x"13",  x"c2",  x"5c",  x"e1",  x"94",  x"72",  x"f3",  x"c1", -- 0F38
         x"22",  x"f2",  x"28",  x"23",  x"88",  x"af",  x"c6",  x"0c", -- 0F40
         x"92",  x"d3",  x"58",  x"ff",  x"c0",  x"58",  x"8c",  x"c9", -- 0F48
         x"75",  x"31",  x"d6",  x"78",  x"b6",  x"b3",  x"76",  x"b2", -- 0F50
         x"a2",  x"2e",  x"14",  x"03",  x"c3",  x"cd",  x"a8",  x"6d", -- 0F58
         x"f2",  x"94",  x"06",  x"c2",  x"bc",  x"98",  x"d4",  x"cd", -- 0F60
         x"07",  x"da",  x"8d",  x"04",  x"0c",  x"d7",  x"92",  x"04", -- 0F68
         x"aa",  x"29",  x"72",  x"7e",  x"82",  x"84",  x"d4",  x"46", -- 0F70
         x"08",  x"dd",  x"33",  x"25",  x"46",  x"fb",  x"b5",  x"0a", -- 0F78
         x"6c",  x"95",  x"46",  x"b2",  x"da",  x"91",  x"19",  x"85", -- 0F80
         x"ce",  x"04",  x"62",  x"ce",  x"66",  x"aa",  x"4a",  x"c8", -- 0F88
         x"11",  x"f3",  x"9c",  x"da",  x"cf",  x"4d",  x"5a",  x"ab", -- 0F90
         x"31",  x"f8",  x"11",  x"05",  x"57",  x"f9",  x"86",  x"3c", -- 0F98
         x"cb",  x"04",  x"03",  x"f8",  x"1e",  x"a3",  x"85",  x"f1", -- 0FA0
         x"31",  x"f9",  x"6c",  x"6e",  x"81",  x"2b",  x"dc",  x"d5", -- 0FA8
         x"a6",  x"f8",  x"d3",  x"c1",  x"04",  x"76",  x"f9",  x"cb", -- 0FB0
         x"70",  x"ad",  x"d3",  x"2c",  x"99",  x"92",  x"89",  x"7d", -- 0FB8
         x"ce",  x"0d",  x"b9",  x"3e",  x"00",  x"98",  x"02",  x"9b", -- 0FC0
         x"9e",  x"02",  x"9a",  x"38",  x"a7",  x"8a",  x"01",  x"18", -- 0FC8
         x"66",  x"e1",  x"24",  x"e5",  x"84",  x"d7",  x"f4",  x"90", -- 0FD0
         x"d7",  x"9d",  x"f5",  x"05",  x"03",  x"91",  x"f6",  x"05", -- 0FD8
         x"54",  x"09",  x"c5",  x"e6",  x"a9",  x"96",  x"66",  x"f4", -- 0FE0
         x"a8",  x"9e",  x"33",  x"f5",  x"7b",  x"03",  x"f6",  x"7a", -- 0FE8
         x"03",  x"79",  x"f7",  x"31",  x"7a",  x"18",  x"34",  x"28", -- 0FF0
         x"a5",  x"4c",  x"c3",  x"39",  x"95",  x"48",  x"e3",  x"24", -- 0FF8
         x"45",  x"4c",  x"a1",  x"d8",  x"ae",  x"13",  x"71",  x"15", -- 1000
         x"51",  x"b5",  x"a0",  x"a2",  x"ce",  x"c3",  x"81",  x"a1", -- 1008
         x"77",  x"8c",  x"e8",  x"79",  x"e9",  x"ce",  x"a0",  x"a5", -- 1010
         x"68",  x"96",  x"68",  x"db",  x"c2",  x"a7",  x"99",  x"8d", -- 1018
         x"ae",  x"c4",  x"fe",  x"a3",  x"da",  x"20",  x"d8",  x"dd", -- 1020
         x"48",  x"03",  x"fe",  x"7a",  x"c7",  x"15",  x"6f",  x"bd", -- 1028
         x"d6",  x"25",  x"00",  x"e3",  x"6a",  x"66",  x"11",  x"81", -- 1030
         x"19",  x"98",  x"aa",  x"44",  x"21",  x"20",  x"00",  x"e5", -- 1038
         x"f1",  x"84",  x"e9",  x"cd",  x"82",  x"19",  x"b0",  x"3f", -- 1040
         x"92",  x"b0",  x"16",  x"ea",  x"76",  x"02",  x"b9",  x"7a", -- 1048
         x"d1",  x"a6",  x"4e",  x"2b",  x"1f",  x"7e",  x"09",  x"f0", -- 1050
         x"13",  x"cc",  x"19",  x"40",  x"01",  x"0b",  x"c7",  x"d7", -- 1058
         x"96",  x"a5",  x"27",  x"68",  x"5d",  x"23",  x"4d",  x"24", -- 1060
         x"f4",  x"aa",  x"23",  x"d5",  x"1c",  x"eb",  x"0c",  x"92", -- 1068
         x"98",  x"34",  x"bb",  x"ef",  x"00",  x"d1",  x"94",  x"89", -- 1070
         x"28",  x"11",  x"70",  x"26",  x"11",  x"69",  x"97",  x"f1", -- 1078
         x"55",  x"c2",  x"4c",  x"ca",  x"05",  x"99",  x"6a",  x"3c", -- 1080
         x"d9",  x"15",  x"3b",  x"f6",  x"68",  x"03",  x"e0",  x"ce", -- 1088
         x"84",  x"8e",  x"ab",  x"64",  x"8f",  x"f8",  x"f4",  x"b0", -- 1090
         x"b1",  x"12",  x"ca",  x"6d",  x"9a",  x"d4",  x"56",  x"c3", -- 1098
         x"c4",  x"86",  x"e5",  x"dc",  x"98",  x"cf",  x"11",  x"74", -- 10A0
         x"fb",  x"41",  x"d9",  x"8c",  x"e9",  x"2a",  x"d9",  x"0a", -- 10A8
         x"3e",  x"d9",  x"05",  x"3e",  x"30",  x"58",  x"f9",  x"d1", -- 10B0
         x"4b",  x"39",  x"21",  x"db",  x"55",  x"8d",  x"50",  x"86", -- 10B8
         x"16",  x"18",  x"28",  x"de",  x"00",  x"7e",  x"e6",  x"3f", -- 10C0
         x"67",  x"7a",  x"03",  x"fe",  x"e5",  x"28",  x"08",  x"d6", -- 10C8
         x"2e",  x"2d",  x"08",  x"cb",  x"5c",  x"28",  x"13",  x"a0", -- 10D0
         x"c4",  x"ef",  x"65",  x"ce",  x"14",  x"d8",  x"ff",  x"39", -- 10D8
         x"3e",  x"28",  x"0f",  x"28",  x"9a",  x"5b",  x"f8",  x"2f", -- 10E0
         x"23",  x"04",  x"0e",  x"47",  x"f9",  x"02",  x"dd",  x"3b", -- 10E8
         x"52",  x"b7",  x"a6",  x"da",  x"a4",  x"ad",  x"be",  x"04", -- 10F0
         x"cf",  x"16",  x"e5",  x"a4",  x"27",  x"01",  x"20",  x"03", -- 10F8
         x"ac",  x"4f",  x"0f",  x"a6",  x"77",  x"77",  x"fd",  x"2a", -- 1100
         x"be",  x"f3",  x"c4",  x"7c",  x"93",  x"ee",  x"c6",  x"07", -- 1108
         x"b7",  x"c0",  x"61",  x"5e",  x"aa",  x"c6",  x"aa",  x"b9", -- 1110
         x"c3",  x"60",  x"04",  x"6c",  x"da",  x"00",  x"19",  x"4e", -- 1118
         x"3e",  x"20",  x"60",  x"91",  x"ad",  x"17",  x"a1",  x"97", -- 1120
         x"c0",  x"6f",  x"42",  x"79",  x"fe",  x"2f",  x"28",  x"3d", -- 1128
         x"c1",  x"95",  x"20",  x"60",  x"c3",  x"01",  x"30",  x"af", -- 1130
         x"67",  x"b5",  x"5b",  x"08",  x"cc",  x"05",  x"96",  x"fe", -- 1138
         x"38",  x"14",  x"08",  x"b4",  x"d6",  x"08",  x"20",  x"0a", -- 1140
         x"21",  x"b4",  x"28",  x"1e",  x"4f",  x"f1",  x"15",  x"4f", -- 1148
         x"0b",  x"18",  x"bf",  x"e6",  x"78",  x"1b",  x"34",  x"fd", -- 1150
         x"d1",  x"83",  x"86",  x"fb",  x"6f",  x"41",  x"f4",  x"ad", -- 1158
         x"fc",  x"67",  x"0a",  x"71",  x"18",  x"ab",  x"68",  x"52", -- 1160
         x"32",  x"fd",  x"75",  x"60",  x"74",  x"01",  x"9c",  x"e4", -- 1168
         x"c6",  x"0b",  x"a7",  x"d1",  x"48",  x"fc",  x"d1",  x"ef", -- 1170
         x"ff",  x"d1",  x"ea",  x"65",  x"20",  x"9d",  x"50",  x"12", -- 1178
         x"82",  x"81",  x"7d",  x"22",  x"55",  x"92",  x"a1",  x"09", -- 1180
         x"62",  x"a1",  x"46",  x"09",  x"15",  x"a1",  x"85",  x"e4", -- 1188
         x"9c",  x"df",  x"a4",  x"a5",  x"7e",  x"b2",  x"a4",  x"02", -- 1190
         x"5c",  x"9c",  x"c1",  x"c5",  x"1e",  x"00",  x"51",  x"e0", -- 1198
         x"53",  x"16",  x"91",  x"62",  x"d1",  x"20",  x"c4",  x"b0", -- 11A0
         x"d6",  x"05",  x"66",  x"20",  x"d5",  x"e5",  x"06",  x"7a", -- 11A8
         x"02",  x"03",  x"1c",  x"7b",  x"ae",  x"01",  x"38",  x"e2", -- 11B0
         x"33",  x"33",  x"31",  x"a3",  x"1f",  x"11",  x"08",  x"21", -- 11B8
         x"c6",  x"18",  x"20",  x"1f",  x"3e",  x"2e",  x"dc",  x"1b", -- 11C0
         x"1e",  x"69",  x"fe",  x"35",  x"68",  x"13",  x"08",  x"90", -- 11C8
         x"2d",  x"0b",  x"38",  x"5d",  x"ea",  x"2d",  x"bd",  x"80", -- 11D0
         x"d5",  x"f8",  x"84",  x"b4",  x"92",  x"24",  x"15",  x"b0", -- 11D8
         x"48",  x"d6",  x"06",  x"c6",  x"1c",  x"5e",  x"6f",  x"99", -- 11E0
         x"75",  x"c9",  x"6f",  x"d5",  x"82",  x"85",  x"4e",  x"52", -- 11E8
         x"b4",  x"b7",  x"b8",  x"a5",  x"e3",  x"b7",  x"37",  x"04", -- 11F0
         x"31",  x"6b",  x"37",  x"5f",  x"2b",  x"4d",  x"18",  x"2b", -- 11F8
         x"44",  x"27",  x"6a",  x"63",  x"c8",  x"1f",  x"06",  x"a4", -- 1200
         x"1f",  x"16",  x"76",  x"1f",  x"b5",  x"48",  x"36",  x"e8", -- 1208
         x"fb",  x"54",  x"f6",  x"fb",  x"6c",  x"62",  x"08",  x"62", -- 1210
         x"09",  x"46",  x"f0",  x"d4",  x"13",  x"78",  x"c0",  x"bb", -- 1218
         x"20",  x"0a",  x"f3",  x"d8",  x"f2",  x"8c",  x"10",  x"72", -- 1220
         x"09",  x"33",  x"18",  x"ed",  x"a5",  x"cd",  x"07",  x"74", -- 1228
         x"09",  x"14",  x"2f",  x"9c",  x"d6",  x"b2",  x"12",  x"df", -- 1230
         x"a3",  x"a0",  x"d3",  x"d4",  x"83",  x"a1",  x"9c",  x"14", -- 1238
         x"b8",  x"77",  x"48",  x"42",  x"80",  x"30",  x"2d",  x"11", -- 1240
         x"c5",  x"e2",  x"92",  x"55",  x"86",  x"db",  x"73",  x"c3", -- 1248
         x"0c",  x"61",  x"9d",  x"dd",  x"71",  x"e7",  x"55",  x"70", -- 1250
         x"bd",  x"6b",  x"06",  x"f7",  x"8b",  x"f1",  x"7d",  x"e3", -- 1258
         x"3d",  x"91",  x"67",  x"39",  x"bd",  x"99",  x"28",  x"8a", -- 1260
         x"9a",  x"bd",  x"a9",  x"c1",  x"d5",  x"49",  x"20",  x"66", -- 1268
         x"d3",  x"e9",  x"13",  x"26",  x"d2",  x"98",  x"13",  x"4a", -- 1270
         x"52",  x"9b",  x"99",  x"f9",  x"df",  x"e8",  x"ac",  x"c5", -- 1278
         x"a5",  x"54",  x"c1",  x"c2",  x"c9",  x"3c",  x"55",  x"9b", -- 1280
         x"11",  x"89",  x"0e",  x"19",  x"cb",  x"66",  x"19",  x"d0", -- 1288
         x"2a",  x"10",  x"a5",  x"a5",  x"fb",  x"95",  x"6e",  x"f8", -- 1290
         x"d3",  x"0e",  x"73",  x"a3",  x"4c",  x"74",  x"f7",  x"a5", -- 1298
         x"06",  x"f6",  x"dd",  x"5e",  x"a2",  x"01",  x"56",  x"ff", -- 12A0
         x"21",  x"02",  x"3d",  x"c1",  x"91",  x"18",  x"88",  x"ad", -- 12A8
         x"ba",  x"40",  x"19",  x"e5",  x"21",  x"fe",  x"01",  x"e5", -- 12B0
         x"94",  x"bb",  x"11",  x"e5",  x"dd",  x"c8",  x"18",  x"f2", -- 12B8
         x"b7",  x"db",  x"47",  x"3a",  x"9e",  x"4d",  x"98",  x"1a", -- 12C0
         x"5e",  x"05",  x"ce",  x"e2",  x"d3",  x"66",  x"c5",  x"99", -- 12C8
         x"55",  x"d0",  x"f0",  x"7c",  x"d6",  x"aa",  x"a5",  x"19", -- 12D0
         x"02",  x"2c",  x"19",  x"d5",  x"4b",  x"2e",  x"36",  x"82", -- 12D8
         x"16",  x"4a",  x"d1",  x"c1",  x"09",  x"12",  x"9a",  x"40", -- 12E0
         x"46",  x"fb",  x"60",  x"40",  x"41",  x"20",  x"03",  x"6f", -- 12E8
         x"18",  x"4a",  x"41",  x"3e",  x"52",  x"82",  x"7b",  x"3e", -- 12F0
         x"9c",  x"98",  x"a7",  x"3e",  x"02",  x"d4",  x"51",  x"60", -- 12F8
         x"d5",  x"be",  x"a2",  x"d7",  x"dd",  x"c4",  x"b2",  x"89", -- 1300
         x"fa",  x"21",  x"21",  x"40",  x"04",  x"cd",  x"9a",  x"8f", -- 1308
         x"7d",  x"0f",  x"58",  x"30",  x"a5",  x"0c",  x"7c",  x"a2", -- 1310
         x"af",  x"fa",  x"5b",  x"c2",  x"02",  x"c3",  x"02",  x"6a", -- 1318
         x"c4",  x"02",  x"c5",  x"e0",  x"d4",  x"39",  x"a4",  x"ca", -- 1320
         x"eb",  x"fb",  x"37",  x"7d",  x"03",  x"ec",  x"b2",  x"67", -- 1328
         x"9d",  x"a6",  x"cf",  x"48",  x"55",  x"eb",  x"71",  x"4a", -- 1330
         x"9d",  x"7a",  x"ed",  x"e3",  x"68",  x"96",  x"ff",  x"2a", -- 1338
         x"46",  x"60",  x"ff",  x"a8",  x"10",  x"fc",  x"26",  x"61", -- 1340
         x"b3",  x"67",  x"32",  x"46",  x"c5",  x"82",  x"9d",  x"28", -- 1348
         x"c9",  x"90",  x"3c",  x"29",  x"b8",  x"34",  x"7e",  x"0d", -- 1350
         x"32",  x"5a",  x"ed",  x"67",  x"bb",  x"3f",  x"dd",  x"4a", -- 1358
         x"98",  x"5b",  x"25",  x"c4",  x"25",  x"cf",  x"85",  x"06", -- 1360
         x"68",  x"c2",  x"06",  x"c3",  x"85",  x"7b",  x"7a",  x"7d", -- 1368
         x"8a",  x"fe",  x"b0",  x"ad",  x"0b",  x"7a",  x"f6",  x"15", -- 1370
         x"06",  x"4c",  x"08",  x"c7",  x"4a",  x"24",  x"a2",  x"12", -- 1378
         x"0d",  x"e5",  x"3e",  x"35",  x"38",  x"a6",  x"ae",  x"38", -- 1380
         x"46",  x"dc",  x"48",  x"6f",  x"74",  x"67",  x"a6",  x"ce", -- 1388
         x"61",  x"11",  x"a6",  x"72",  x"f3",  x"20",  x"5a",  x"13", -- 1390
         x"17",  x"17",  x"78",  x"17",  x"bf",  x"9c",  x"49",  x"23", -- 1398
         x"dd",  x"0a",  x"f8",  x"bf",  x"9a",  x"c7",  x"85",  x"fa", -- 13A0
         x"13",  x"03",  x"fb",  x"00",  x"57",  x"81",  x"06",  x"9e", -- 13A8
         x"15",  x"66",  x"f9",  x"66",  x"e6",  x"05",  x"52",  x"a8", -- 13B0
         x"05",  x"9d",  x"4b",  x"bc",  x"be",  x"b0",  x"1e",  x"96", -- 13B8
         x"0c",  x"73",  x"c0",  x"e7",  x"d2",  x"c1",  x"57",  x"f1", -- 13C0
         x"1e",  x"74",  x"f1",  x"f9",  x"c5",  x"05",  x"f8",  x"c6", -- 13C8
         x"0a",  x"6d",  x"c4",  x"4d",  x"d4",  x"89",  x"b1",  x"f7", -- 13D0
         x"e5",  x"37",  x"58",  x"e7",  x"aa",  x"e1",  x"ec",  x"d5", -- 13D8
         x"e1",  x"59",  x"6d",  x"9b",  x"0a",  x"7e",  x"c2",  x"81", -- 13E0
         x"a1",  x"62",  x"c3",  x"88",  x"84",  x"90",  x"c4",  x"8d", -- 13E8
         x"63",  x"4f",  x"04",  x"c5",  x"8c",  x"47",  x"27",  x"c8", -- 13F0
         x"33",  x"66",  x"f7",  x"8f",  x"9c",  x"d5",  x"45",  x"02", -- 13F8
         x"96",  x"d3",  x"26",  x"45",  x"f5",  x"a3",  x"bf",  x"06", -- 1400
         x"11",  x"17",  x"66",  x"f5",  x"77",  x"1d",  x"49",  x"71", -- 1408
         x"f2",  x"92",  x"1d",  x"f3",  x"8d",  x"e5",  x"3f",  x"ab", -- 1410
         x"08",  x"95",  x"13",  x"66",  x"f3",  x"43",  x"23",  x"83", -- 1418
         x"c6",  x"01",  x"f8",  x"7b",  x"b2",  x"38",  x"f8",  x"22", -- 1420
         x"13",  x"82",  x"f8",  x"8c",  x"33",  x"fd",  x"66",  x"b3", -- 1428
         x"59",  x"6e",  x"b6",  x"98",  x"74",  x"ee",  x"d1",  x"30", -- 1430
         x"ef",  x"ef",  x"50",  x"f0",  x"f3",  x"15",  x"f1",  x"00", -- 1438
         x"fb",  x"c5",  x"ee",  x"6f",  x"73",  x"fc",  x"ef",  x"bb", -- 1440
         x"bc",  x"04",  x"f0",  x"4f",  x"af",  x"82",  x"1b",  x"f1", -- 1448
         x"47",  x"7d",  x"13",  x"be",  x"6b",  x"36",  x"ee",  x"7c", -- 1450
         x"0b",  x"bf",  x"06",  x"ef",  x"cd",  x"21",  x"9e",  x"c0", -- 1458
         x"06",  x"f0",  x"4d",  x"23",  x"c1",  x"06",  x"f1",  x"2e", -- 1460
         x"77",  x"c5",  x"27",  x"66",  x"06",  x"e3",  x"60",  x"3c", -- 1468
         x"cb",  x"1b",  x"10",  x"fa",  x"58",  x"01",  x"e3",  x"15", -- 1470
         x"ee",  x"93",  x"2f",  x"95",  x"06",  x"ef",  x"9c",  x"2f", -- 1478
         x"95",  x"06",  x"f0",  x"99",  x"2f",  x"92",  x"06",  x"f1", -- 1480
         x"98",  x"58",  x"2f",  x"c7",  x"39",  x"5e",  x"94",  x"90", -- 1488
         x"eb",  x"fc",  x"0d",  x"17",  x"66",  x"f1",  x"a1",  x"a8", -- 1490
         x"cd",  x"2c",  x"66",  x"ef",  x"e4",  x"12",  x"5e",  x"0b", -- 1498
         x"df",  x"7d",  x"ff",  x"02",  x"6f",  x"7c",  x"81",  x"a5", -- 14A0
         x"7b",  x"50",  x"c5",  x"7a",  x"a3",  x"b3",  x"c9",  x"db", -- 14A8
         x"06",  x"b1",  x"52",  x"4e",  x"e4",  x"09",  x"46",  x"f9", -- 14B0
         x"fd",  x"09",  x"68",  x"f4",  x"fd",  x"73",  x"0c",  x"02", -- 14B8
         x"fd",  x"72",  x"03",  x"15",  x"7d",  x"d6",  x"03",  x"f7", -- 14C0
         x"7c",  x"de",  x"0f",  x"7b",  x"de",  x"db",  x"2c",  x"02", -- 14C8
         x"30",  x"02",  x"24",  x"06",  x"01",  x"0f",  x"4b",  x"ff", -- 14D0
         x"0f",  x"56",  x"87",  x"4f",  x"d1",  x"0f",  x"f8",  x"03", -- 14D8
         x"1f",  x"38",  x"06",  x"79",  x"9b",  x"3d",  x"23",  x"02", -- 14E0
         x"b3",  x"05",  x"20",  x"05",  x"03",  x"78",  x"05",  x"98", -- 14E8
         x"d7",  x"e4",  x"dc",  x"29",  x"05",  x"f5",  x"0e",  x"61", -- 14F0
         x"b3",  x"28",  x"d7",  x"94",  x"ef",  x"78",  x"81",  x"8b", -- 14F8
         x"31",  x"b2",  x"14",  x"1f",  x"84",  x"8a",  x"ff",  x"94", -- 1500
         x"8a",  x"98",  x"5e",  x"0a",  x"56",  x"f5",  x"21",  x"44", -- 1508
         x"2c",  x"a6",  x"c2",  x"2f",  x"56",  x"5c",  x"ef",  x"0f", -- 1510
         x"86",  x"0e",  x"18",  x"43",  x"10",  x"f6",  x"d1",  x"10", -- 1518
         x"f7",  x"47",  x"20",  x"7e",  x"ea",  x"b6",  x"94",  x"ba", -- 1520
         x"39",  x"05",  x"7e",  x"eb",  x"e5",  x"b9",  x"0e",  x"bc", -- 1528
         x"05",  x"7e",  x"74",  x"ec",  x"08",  x"be",  x"39",  x"05", -- 1530
         x"7e",  x"ed",  x"d0",  x"08",  x"c0",  x"a3",  x"ed",  x"95", -- 1538
         x"44",  x"fd",  x"96",  x"3b",  x"12",  x"f8",  x"12",  x"c1", -- 1540
         x"ec",  x"19",  x"29",  x"97",  x"cb",  x"88",  x"7b",  x"ec", -- 1548
         x"4a",  x"49",  x"7b",  x"95",  x"47",  x"78",  x"2a",  x"45", -- 1550
         x"7c",  x"69",  x"43",  x"89",  x"84",  x"56",  x"44",  x"84", -- 1558
         x"3a",  x"b2",  x"84",  x"b3",  x"e8",  x"ca",  x"7b",  x"83", -- 1560
         x"5f",  x"77",  x"28",  x"8a",  x"57",  x"73",  x"8c",  x"67", -- 1568
         x"a3",  x"6f",  x"8d",  x"6f",  x"b7",  x"1c",  x"bd",  x"58", -- 1570
         x"72",  x"bd",  x"b1",  x"74",  x"bd",  x"25",  x"75",  x"03", -- 1578
         x"f8",  x"06",  x"23",  x"9c",  x"f2",  x"b7",  x"08",  x"22", -- 1580
         x"ac",  x"8e",  x"ac",  x"d2",  x"21",  x"ba",  x"9c",  x"c3", -- 1588
         x"ed",  x"4b",  x"ca",  x"17",  x"78",  x"b1",  x"ab",  x"10", -- 1590
         x"05",  x"c3",  x"73",  x"a3",  x"23",  x"21",  x"01",  x"6b", -- 1598
         x"f8",  x"3b",  x"b0",  x"b6",  x"d8",  x"11",  x"fc",  x"11", -- 15A0
         x"fd",  x"eb",  x"13",  x"6f",  x"13",  x"ef",  x"6d",  x"0c", -- 15A8
         x"fa",  x"0c",  x"fb",  x"94",  x"6c",  x"fa",  x"12",  x"f0", -- 15B0
         x"65",  x"fb",  x"12",  x"62",  x"48",  x"8a",  x"d5",  x"d3", -- 15B8
         x"ff",  x"2c",  x"cf",  x"23",  x"6e",  x"fd",  x"19",  x"1c", -- 15C0
         x"09",  x"75",  x"fb",  x"c5",  x"d5",  x"a3",  x"d3",  x"93", -- 15C8
         x"59",  x"94",  x"e0",  x"cd",  x"65",  x"51",  x"9c",  x"f6", -- 15D0
         x"1b",  x"d1",  x"c1",  x"bc",  x"0c",  x"20",  x"74",  x"1a", -- 15D8
         x"a4",  x"94",  x"09",  x"30",  x"fd",  x"1b",  x"cb",  x"0b", -- 15E0
         x"66",  x"c7",  x"f2",  x"f0",  x"18",  x"3d",  x"63",  x"21", -- 15E8
         x"fd",  x"bd",  x"10",  x"e4",  x"f8",  x"04",  x"42",  x"dc", -- 15F0
         x"b6",  x"32",  x"e1",  x"95",  x"dc",  x"b9",  x"27",  x"40", -- 15F8
         x"dc",  x"a6",  x"d1",  x"bd",  x"2c",  x"1a",  x"e1",  x"07", -- 1600
         x"09",  x"21",  x"1c",  x"97",  x"76",  x"b5",  x"3b",  x"d0", -- 1608
         x"3b",  x"2b",  x"b4",  x"c3",  x"f0",  x"11",  x"4c",  x"73", -- 1610
         x"f3",  x"07",  x"21",  x"16",  x"4b",  x"15",  x"ad",  x"92", -- 1618
         x"02",  x"c3",  x"01",  x"3c",  x"f6",  x"17",  x"da",  x"92", -- 1620
         x"b6",  x"d6",  x"cb",  x"dc",  x"d6",  x"6d",  x"26",  x"2a", -- 1628
         x"8a",  x"81",  x"e3",  x"33",  x"b6",  x"e2",  x"33",  x"f4", -- 1630
         x"0f",  x"09",  x"db",  x"dd",  x"b6",  x"da",  x"04",  x"9c", -- 1638
         x"21",  x"a7",  x"c5",  x"0c",  x"da",  x"c6",  x"01",  x"cf", -- 1640
         x"af",  x"14",  x"37",  x"cd",  x"c9",  x"ff",  x"06",  x"0f", -- 1648
         x"38",  x"1e",  x"04",  x"ac",  x"1e",  x"c0",  x"09",  x"11", -- 1650
         x"1a",  x"fd",  x"d8",  x"56",  x"6b",  x"2b",  x"16",  x"88", -- 1658
         x"d9",  x"58",  x"2b",  x"fb",  x"c4",  x"65",  x"f2",  x"96", -- 1660
         x"0c",  x"56",  x"fb",  x"c1",  x"29",  x"eb",  x"82",  x"ca", -- 1668
         x"98",  x"88",  x"f6",  x"4f",  x"a5",  x"e4",  x"29",  x"f7", -- 1670
         x"47",  x"83",  x"9a",  x"f8",  x"88",  x"e4",  x"04",  x"f9", -- 1678
         x"67",  x"9a",  x"be",  x"f6",  x"93",  x"be",  x"70",  x"fe", -- 1680
         x"17",  x"36",  x"f8",  x"00",  x"ac",  x"17",  x"27",  x"76", -- 1688
         x"26",  x"25",  x"7c",  x"a6",  x"24",  x"30",  x"22",  x"71", -- 1690
         x"cb",  x"02",  x"70",  x"07",  x"63",  x"5c",  x"22",  x"2d", -- 1698
         x"bf",  x"63",  x"2f",  x"0f",  x"69",  x"ca",  x"da",  x"0d", -- 16A0
         x"c8",  x"5a",  x"0b",  x"f2",  x"45",  x"0b",  x"f3",  x"ad", -- 16A8
         x"27",  x"26",  x"9f",  x"a5",  x"27",  x"58",  x"f1",  x"f4", -- 16B0
         x"05",  x"b6",  x"04",  x"d6",  x"01",  x"2d",  x"bf",  x"b7", -- 16B8
         x"bc",  x"6b",  x"84",  x"0d",  x"06",  x"ca",  x"1f",  x"a7", -- 16C0
         x"c0",  x"a0",  x"11",  x"89",  x"da",  x"40",  x"eb",  x"b7", -- 16C8
         x"c2",  x"f8",  x"05",  x"a5",  x"dd",  x"cb",  x"ec",  x"46", -- 16D0
         x"52",  x"06",  x"9a",  x"bd",  x"eb",  x"1e",  x"d4",  x"1a", -- 16D8
         x"4e",  x"8a",  x"00",  x"46",  x"ee",  x"f1",  x"3e",  x"09", -- 16E0
         x"cb",  x"38",  x"7c",  x"cb",  x"99",  x"1a",  x"d3",  x"89", -- 16E8
         x"b3",  x"b4",  x"f5",  x"a9",  x"9b",  x"91",  x"8b",  x"66", -- 16F0
         x"25",  x"93",  x"b3",  x"e7",  x"b0",  x"05",  x"e8",  x"02", -- 16F8
         x"b4",  x"e9",  x"9c",  x"03",  x"ea",  x"96",  x"0d",  x"dd", -- 1700
         x"a6",  x"e7",  x"e4",  x"f3",  x"04",  x"e8",  x"79",  x"03", -- 1708
         x"36",  x"e9",  x"78",  x"03",  x"ea",  x"1f",  x"de",  x"6f", -- 1710
         x"7c",  x"53",  x"9e",  x"53",  x"be",  x"7f",  x"73",  x"48", -- 1718
         x"61",  x"b6",  x"4e",  x"b6",  x"eb",  x"20",  x"1f",  x"2b", -- 1720
         x"b0",  x"b3",  x"11",  x"85",  x"55",  x"19",  x"9e",  x"2e", -- 1728
         x"e1",  x"a3",  x"96",  x"e2",  x"04",  x"e3",  x"b1",  x"04", -- 1730
         x"e4",  x"18",  x"3d",  x"32",  x"f2",  x"a7",  x"0d",  x"97", -- 1738
         x"0d",  x"2e",  x"e9",  x"a8",  x"2e",  x"ea",  x"d9",  x"f3", -- 1740
         x"6b",  x"66",  x"e8",  x"b0",  x"32",  x"99",  x"92",  x"a9", -- 1748
         x"af",  x"72",  x"b3",  x"5a",  x"73",  x"15",  x"74",  x"e8", -- 1750
         x"b1",  x"31",  x"e7",  x"21",  x"07",  x"57",  x"28",  x"2d", -- 1758
         x"23",  x"2c",  x"3e",  x"b0",  x"23",  x"be",  x"e1",  x"e8", -- 1760
         x"0c",  x"b5",  x"56",  x"e2",  x"04",  x"e3",  x"b1",  x"04", -- 1768
         x"e4",  x"38",  x"0d",  x"29",  x"b9",  x"69",  x"dc",  x"dd", -- 1770
         x"c7",  x"94",  x"d6",  x"a9",  x"5f",  x"07",  x"a5",  x"31", -- 1778
         x"92",  x"6a",  x"c2",  x"25",  x"23",  x"16",  x"ca",  x"92", -- 1780
         x"83",  x"cd",  x"42",  x"95",  x"5f",  x"ec",  x"d8",  x"b4", -- 1788
         x"b5",  x"47",  x"20",  x"18",  x"35",  x"7e",  x"de",  x"9d", -- 1790
         x"46",  x"07",  x"ed",  x"c3",  x"22",  x"86",  x"e7",  x"47", -- 1798
         x"99",  x"ae",  x"e8",  x"ce",  x"d2",  x"04",  x"e9",  x"cb", -- 17A0
         x"ce",  x"04",  x"25",  x"ea",  x"57",  x"fd",  x"85",  x"70", -- 17A8
         x"57",  x"f5",  x"f9",  x"49",  x"72",  x"56",  x"8b",  x"66", -- 17B0
         x"ec",  x"c0",  x"b2",  x"e7",  x"7b",  x"51",  x"e6",  x"cd", -- 17B8
         x"be",  x"e8",  x"ad",  x"63",  x"96",  x"46",  x"77",  x"df", -- 17C0
         x"3e",  x"91",  x"b3",  x"9e",  x"e8",  x"07",  x"59",  x"e0", -- 17C8
         x"80",  x"96",  x"96",  x"df",  x"94",  x"41",  x"9e",  x"e0", -- 17D0
         x"30",  x"0c",  x"21",  x"8e",  x"dd",  x"0d",  x"b2",  x"19", -- 17D8
         x"5e",  x"4b",  x"56",  x"f1",  x"2c",  x"9f",  x"9a",  x"ef", -- 17E0
         x"c9",  x"b5",  x"0a",  x"79",  x"e5",  x"0a",  x"7d",  x"e6", -- 17E8
         x"00",  x"18",  x"2b",  x"6d",  x"dc",  x"25",  x"e5",  x"05", -- 17F0
         x"dd",  x"bc",  x"05",  x"e6",  x"6a",  x"34",  x"66",  x"e0", -- 17F8
         x"9c",  x"a3",  x"76",  x"06",  x"ed",  x"06",  x"ee",  x"a6", -- 1800
         x"06",  x"eb",  x"06",  x"ec",  x"ac",  x"06",  x"02",  x"66", -- 1808
         x"e6",  x"46",  x"e5",  x"ec",  x"d2",  x"78",  x"92",  x"d9", -- 1810
         x"8a",  x"c5",  x"0b",  x"f2",  x"66",  x"4e",  x"16",  x"6e", -- 1818
         x"e0",  x"11",  x"f2",  x"e5",  x"e7",  x"84",  x"60",  x"d1", -- 1820
         x"e8",  x"8d",  x"47",  x"ca",  x"04",  x"e9",  x"8b",  x"fc", -- 1828
         x"76",  x"ea",  x"fc",  x"f2",  x"85",  x"d6",  x"65",  x"d7", -- 1830
         x"85",  x"e3",  x"83",  x"84",  x"86",  x"2c",  x"b5",  x"d9", -- 1838
         x"c0",  x"87",  x"8e",  x"e0",  x"a5",  x"dc",  x"98",  x"d0", -- 1840
         x"09",  x"77",  x"06",  x"43",  x"d3",  x"08",  x"4a",  x"07", -- 1848
         x"de",  x"ab",  x"56",  x"f0",  x"8c",  x"2a",  x"57",  x"7c", -- 1850
         x"a4",  x"26",  x"5f",  x"b5",  x"12",  x"db",  x"82",  x"c3", -- 1858
         x"8e",  x"a4",  x"3d",  x"ad",  x"94",  x"d1",  x"ad",  x"d4", -- 1860
         x"a1",  x"cc",  x"7c",  x"81",  x"b3",  x"39",  x"36",  x"fd", -- 1868
         x"88",  x"62",  x"c7",  x"a7",  x"46",  x"bb",  x"ed",  x"30", -- 1870
         x"bb",  x"92",  x"ff",  x"fc",  x"b5",  x"b0",  x"9a",  x"45", -- 1878
         x"38",  x"4c",  x"78",  x"94",  x"49",  x"79",  x"92",  x"07", -- 1880
         x"5d",  x"54",  x"83",  x"0c",  x"4e",  x"72",  x"46",  x"07", -- 1888
         x"4d",  x"c5",  x"a3",  x"d3",  x"c6",  x"82",  x"a1",  x"6a", -- 1890
         x"fd",  x"84",  x"85",  x"43",  x"42",  x"84",  x"2b",  x"78", -- 1898
         x"84",  x"5d",  x"1e",  x"85",  x"a6",  x"04",  x"b8",  x"df", -- 18A0
         x"b1",  x"2e",  x"82",  x"04",  x"4d",  x"44",  x"e1",  x"c0", -- 18A8
         x"d0",  x"18",  x"f6",  x"6a",  x"74",  x"03",  x"1b",  x"fd", -- 18B0
         x"d3",  x"34",  x"0e",  x"8a",  x"49",  x"68",  x"96",  x"f1", -- 18B8
         x"46",  x"b8",  x"ee",  x"8c",  x"a8",  x"04",  x"d2",  x"4c", -- 18C0
         x"cd",  x"f0",  x"d7",  x"05",  x"30",  x"18",  x"65",  x"9a", -- 18C8
         x"c0",  x"3b",  x"56",  x"05",  x"4b",  x"42",  x"03",  x"03", -- 18D0
         x"b0",  x"9c",  x"9a",  x"d6",  x"77",  x"6a",  x"02",  x"4d", -- 18D8
         x"a5",  x"69",  x"02",  x"f6",  x"5c",  x"d2",  x"16",  x"d5", -- 18E0
         x"4d",  x"18",  x"58",  x"39",  x"b3",  x"74",  x"7a",  x"7c", -- 18E8
         x"ac",  x"49",  x"99",  x"a7",  x"35",  x"9c",  x"85",  x"01", -- 18F0
         x"6f",  x"03",  x"a8",  x"20",  x"65",  x"6e",  x"06",  x"73", -- 18F8
         x"07",  x"9b",  x"72",  x"19",  x"54",  x"9b",  x"82",  x"bf", -- 1900
         x"69",  x"d8",  x"09",  x"cd",  x"69",  x"97",  x"f1",  x"64", -- 1908
         x"23",  x"82",  x"00",  x"c3",  x"83",  x"ad",  x"c3",  x"00", -- 1910
         x"f5",  x"a9",  x"c3",  x"99",  x"aa",  x"c3",  x"56",  x"ab", -- 1918
         x"00",  x"c3",  x"28",  x"ac",  x"3e",  x"05",  x"cf",  x"c3", -- 1920
         x"0c",  x"90",  x"05",  x"de",  x"a8",  x"b2",  x"05",  x"26", -- 1928
         x"a9",  x"d2",  x"05",  x"e2",  x"24",  x"05",  x"e7",  x"11", -- 1930
         x"48",  x"a3",  x"0b",  x"bc",  x"91",  x"05",  x"2e",  x"22", -- 1938
         x"05",  x"c7",  x"44",  x"17",  x"ce",  x"89",  x"0b",  x"88", -- 1940
         x"12",  x"05",  x"67",  x"24",  x"05",  x"d8",  x"05",  x"48", -- 1948
         x"94",  x"05",  x"76",  x"91",  x"05",  x"b0",  x"20",  x"05", -- 1950
         x"d3",  x"a8",  x"21",  x"60",  x"03",  x"b2",  x"5e",  x"00", -- 1958
         x"2b",  x"6e",  x"cd",  x"35",  x"a9",  x"eb",  x"c9",  x"f1", -- 1960
         x"30",  x"e1",  x"d1",  x"bc",  x"11",  x"f5",  x"cd",  x"38", -- 1968
         x"04",  x"0a",  x"c3",  x"f6",  x"e3",  x"1f",  x"7d",  x"07", -- 1970
         x"9f",  x"e7",  x"ef",  x"03",  x"e7",  x"20",  x"aa",  x"17", -- 1978
         x"7c",  x"f5",  x"70",  x"17",  x"bb",  x"97",  x"00",  x"95", -- 1980
         x"6f",  x"9f",  x"94",  x"67",  x"cb",  x"7a",  x"28",  x"c1", -- 1988
         x"09",  x"93",  x"5f",  x"9f",  x"92",  x"57",  x"42",  x"34", -- 1990
         x"f1",  x"d0",  x"47",  x"50",  x"15",  x"78",  x"c9",  x"17", -- 1998
         x"eb",  x"4b",  x"d0",  x"0a",  x"31",  x"47",  x"18",  x"0a", -- 19A0
         x"30",  x"46",  x"26",  x"00",  x"54",  x"d4",  x"af",  x"80", -- 19A8
         x"b2",  x"00",  x"20",  x"10",  x"06",  x"10",  x"ed",  x"6a", -- 19B0
         x"17",  x"93",  x"0c",  x"30",  x"01",  x"83",  x"3f",  x"07", -- 19B8
         x"10",  x"f6",  x"03",  x"5f",  x"c9",  x"06",  x"09",  x"7d", -- 19C0
         x"6c",  x"1c",  x"33",  x"cb",  x"1d",  x"0d",  x"ed",  x"52", -- 19C8
         x"15",  x"00",  x"19",  x"3f",  x"17",  x"10",  x"f5",  x"cb", -- 19D0
         x"10",  x"50",  x"61",  x"5f",  x"88",  x"10",  x"38",  x"cd", -- 19D8
         x"07",  x"f2",  x"a8",  x"c3",  x"1c",  x"a9",  x"0e",  x"ce", -- 19E0
         x"41",  x"8f",  x"04",  x"cd",  x"f6",  x"d2",  x"11",  x"b8", -- 19E8
         x"20",  x"c3",  x"20",  x"b8",  x"1d",  x"90",  x"bb",  x"2e", -- 19F0
         x"cd",  x"ee",  x"27",  x"60",  x"dc",  x"45",  x"f6",  x"02", -- 19F8
         x"45",  x"66",  x"6a",  x"06",  x"08",  x"29",  x"be",  x"6d", -- 1A00
         x"87",  x"b5",  x"66",  x"44",  x"02",  x"11",  x"4e",  x"18", -- 1A08
         x"16",  x"21",  x"02",  x"da",  x"09",  x"23",  x"09",  x"0c", -- 1A10
         x"60",  x"3e",  x"4d",  x"7d",  x"17",  x"9f",  x"eb",  x"db", -- 1A18
         x"03",  x"09",  x"57",  x"c3",  x"14",  x"ac",  x"cc",  x"a5", -- 1A20
         x"f5",  x"f5",  x"51",  x"3b",  x"fa",  x"2d",  x"07",  x"fa", -- 1A28
         x"9a",  x"fb",  x"83",  x"29",  x"19",  x"fd",  x"b3",  x"f9", -- 1A30
         x"b8",  x"95",  x"2c",  x"05",  x"67",  x"05",  x"06",  x"5f", -- 1A38
         x"b3",  x"05",  x"07",  x"57",  x"42",  x"94",  x"e8",  x"b3", -- 1A40
         x"c2",  x"c8",  x"fd",  x"56",  x"07",  x"97",  x"ff",  x"78", -- 1A48
         x"e1",  x"cd",  x"c0",  x"72",  x"9e",  x"c0",  x"b1",  x"89", -- 1A50
         x"7e",  x"0b",  x"36",  x"08",  x"4f",  x"2a",  x"2d",  x"09", -- 1A58
         x"47",  x"05",  x"0a",  x"21",  x"42",  x"0b",  x"67",  x"4f", -- 1A60
         x"36",  x"4e",  x"c6",  x"0d",  x"46",  x"09",  x"3c",  x"0a", -- 1A68
         x"b3",  x"3c",  x"0b",  x"b4",  x"99",  x"b0",  x"25",  x"db", -- 1A70
         x"6c",  x"b4",  x"c5",  x"58",  x"a8",  x"f1",  x"74",  x"00", -- 1A78
         x"7e",  x"78",  x"0f",  x"29",  x"af",  x"95",  x"33",  x"9c", -- 1A80
         x"4a",  x"74",  x"9b",  x"72",  x"23",  x"9a",  x"57",  x"12", -- 1A88
         x"c9",  x"46",  x"e8",  x"28",  x"0b",  x"cb",  x"a4",  x"06", -- 1A90
         x"20",  x"44",  x"f5",  x"2f",  x"cb",  x"33",  x"08",  x"26", -- 1A98
         x"03",  x"09",  x"16",  x"03",  x"7a",  x"0a",  x"03",  x"7d", -- 1AA0
         x"16",  x"d7",  x"fd",  x"7d",  x"b5",  x"fd",  x"ed",  x"7d", -- 1AA8
         x"dc",  x"bb",  x"7d",  x"cb",  x"4c",  x"7d",  x"30",  x"14", -- 1AB0
         x"b2",  x"2b",  x"0b",  x"3e",  x"95",  x"27",  x"1e",  x"2f", -- 1AB8
         x"ed",  x"03",  x"37",  x"1e",  x"bd",  x"42",  x"1c",  x"53", -- 1AC0
         x"18",  x"b3",  x"17",  x"31",  x"26",  x"38",  x"24",  x"19", -- 1AC8
         x"26",  x"77",  x"04",  x"1c",  x"26",  x"77",  x"05",  x"1f", -- 1AD0
         x"99",  x"ae",  x"d4",  x"0b",  x"ae",  x"f0",  x"89",  x"55", -- 1AD8
         x"62",  x"15",  x"d9",  x"c5",  x"20",  x"aa",  x"18",  x"a1", -- 1AE0
         x"31",  x"4c",  x"86",  x"fa",  x"be",  x"dd",  x"98",  x"e2", -- 1AE8
         x"53",  x"ff",  x"0c",  x"e2",  x"82",  x"ab",  x"05",  x"47", -- 1AF0
         x"47",  x"0b",  x"e2",  x"4e",  x"40",  x"4f",  x"46",  x"40", -- 1AF8
         x"84",  x"ef",  x"8d",  x"30",  x"fe",  x"30",  x"21",  x"63", -- 1B00
         x"dc",  x"5d",  x"ba",  x"20",  x"de",  x"d1",  x"a5",  x"48", -- 1B08
         x"e0",  x"35",  x"f6",  x"d2",  x"0d",  x"e2",  x"71",  x"f6", -- 1B10
         x"18",  x"18",  x"df",  x"2c",  x"1f",  x"05",  x"7d",  x"1d", -- 1B18
         x"05",  x"f7",  x"1b",  x"05",  x"19",  x"30",  x"e7",  x"cb", -- 1B20
         x"90",  x"3b",  x"cb",  x"09",  x"c5",  x"cd",  x"5e",  x"87", -- 1B28
         x"f0",  x"b5",  x"22",  x"ae",  x"fe",  x"15",  x"f2",  x"19", -- 1B30
         x"4c",  x"db",  x"44",  x"4d",  x"1a",  x"af",  x"6f",  x"b0", -- 1B38
         x"d8",  x"6f",  x"b6",  x"98",  x"d5",  x"79",  x"29",  x"cb", -- 1B40
         x"2c",  x"11",  x"17",  x"d9",  x"d1",  x"f7",  x"00",  x"d1", -- 1B48
         x"3b",  x"76",  x"01",  x"05",  x"92",  x"42",  x"36",  x"ff", -- 1B50
         x"20",  x"82",  x"d7",  x"c9",  x"96",  x"67",  x"62",  x"93", -- 1B58
         x"04",  x"a2",  x"95",  x"51",  x"05",  x"91",  x"3c",  x"06", -- 1B60
         x"03",  x"13",  x"16",  x"cb",  x"60",  x"20",  x"37",  x"cb", -- 1B68
         x"13",  x"cb",  x"12",  x"cb",  x"07",  x"44",  x"28",  x"02", -- 1B70
         x"cb",  x"c0",  x"ec",  x"ae",  x"96",  x"49",  x"82",  x"be", -- 1B78
         x"bc",  x"b2",  x"0a",  x"7a",  x"b1",  x"e9",  x"5a",  x"18", -- 1B80
         x"11",  x"47",  x"d6",  x"12",  x"4f",  x"13",  x"5f",  x"b5", -- 1B88
         x"14",  x"57",  x"0a",  x"43",  x"c6",  x"dd",  x"35",  x"93", -- 1B90
         x"8c",  x"a6",  x"48",  x"20",  x"a5",  x"b1",  x"ce",  x"45", -- 1B98
         x"33",  x"0e",  x"cf",  x"b0",  x"96",  x"e8",  x"01",  x"b6", -- 1BA0
         x"08",  x"20",  x"05",  x"44",  x"0e",  x"18",  x"5c",  x"68", -- 1BA8
         x"b4",  x"ae",  x"08",  x"87",  x"ac",  x"87",  x"52",  x"ff", -- 1BB0
         x"9a",  x"ea",  x"2b",  x"58",  x"e5",  x"a1",  x"92",  x"2c", -- 1BB8
         x"fd",  x"1a",  x"96",  x"7f",  x"59",  x"39",  x"f9",  x"05", -- 1BC0
         x"12",  x"c9",  x"be",  x"28",  x"0c",  x"58",  x"05",  x"84", -- 1BC8
         x"30",  x"fc",  x"e4",  x"0b",  x"03",  x"13",  x"18",  x"d1", -- 1BD0
         x"bc",  x"9f",  x"0e",  x"9a",  x"57",  x"67",  x"49",  x"4a", -- 1BD8
         x"25",  x"fc",  x"a3",  x"56",  x"bf",  x"be",  x"d1",  x"89", -- 1BE0
         x"84",  x"30",  x"8f",  x"48",  x"cf",  x"80",  x"51",  x"58", -- 1BE8
         x"0b",  x"7b",  x"b2",  x"50",  x"28",  x"6f",  x"06",  x"77", -- 1BF0
         x"23",  x"26",  x"18",  x"f2",  x"19",  x"8a",  x"2a",  x"90", -- 1BF8
         x"93",  x"1f",  x"0a",  x"62",  x"e9",  x"24",  x"18",  x"f9", -- 1C00
         x"a0",  x"9a",  x"1a",  x"73",  x"13",  x"e6",  x"87",  x"d4", -- 1C08
         x"0c",  x"39",  x"2a",  x"c1",  x"e1",  x"a8",  x"8d",  x"af", -- 1C10
         x"47",  x"4f",  x"01",  x"ed",  x"b1",  x"21",  x"ff",  x"ff", -- 1C18
         x"ed",  x"42",  x"1a",  x"ac",  x"75",  x"85",  x"ae",  x"39", -- 1C20
         x"f0",  x"89",  x"23",  x"23",  x"40",  x"bb",  x"69",  x"60", -- 1C28
         x"eb",  x"09",  x"fd",  x"8e",  x"21",  x"0e",  x"14",  x"65", -- 1C30
         x"f7",  x"90",  x"d5",  x"9e",  x"7e",  x"ae",  x"15",  x"6f", -- 1C38
         x"c5",  x"9f",  x"5c",  x"d7",  x"e4",  x"d0",  x"55",  x"22", -- 1C40
         x"5c",  x"c1",  x"33",  x"b0",  x"2e",  x"8b",  x"38",  x"51", -- 1C48
         x"7e",  x"97",  x"d9",  x"04",  x"fb",  x"d1",  x"a4",  x"6f", -- 1C50
         x"d5",  x"47",  x"e2",  x"15",  x"f0",  x"39",  x"37",  x"7e", -- 1C58
         x"fa",  x"85",  x"57",  x"a6",  x"81",  x"23",  x"8c",  x"5f", -- 1C60
         x"13",  x"41",  x"e3",  x"76",  x"75",  x"06",  x"3d",  x"fe", -- 1C68
         x"97",  x"72",  x"37",  x"ce",  x"c2",  x"b3",  x"de",  x"8f", -- 1C70
         x"d4",  x"55",  x"ee",  x"ec",  x"c1",  x"1d",  x"d1",  x"19", -- 1C78
         x"eb",  x"58",  x"65",  x"95",  x"bd",  x"5e",  x"5e",  x"2c", -- 1C80
         x"21",  x"c5",  x"16",  x"1d",  x"eb",  x"99",  x"37",  x"e5", -- 1C88
         x"e7",  x"d8",  x"1b",  x"61",  x"8a",  x"33",  x"0f",  x"7e", -- 1C90
         x"47",  x"c8",  x"6e",  x"66",  x"fa",  x"c3",  x"48",  x"fd", -- 1C98
         x"75",  x"fa",  x"e2",  x"74",  x"01",  x"6a",  x"20",  x"80", -- 1CA0
         x"08",  x"99",  x"3a",  x"e8",  x"34",  x"b6",  x"12",  x"19", -- 1CA8
         x"d1",  x"25",  x"9a",  x"68",  x"b0",  x"17",  x"c1",  x"72", -- 1CB0
         x"77",  x"59",  x"50",  x"0a",  x"4f",  x"2e",  x"1e",  x"9a", -- 1CB8
         x"08",  x"59",  x"a6",  x"4e",  x"d1",  x"be",  x"3e",  x"f6", -- 1CC0
         x"bd",  x"13",  x"fc",  x"b1",  x"e5",  x"fe",  x"c2",  x"d8", -- 1CC8
         x"d4",  x"86",  x"08",  x"5b",  x"6f",  x"d2",  x"0b",  x"8e", -- 1CD0
         x"09",  x"67",  x"d0",  x"66",  x"8e",  x"f0",  x"76",  x"ce", -- 1CD8
         x"c4",  x"8e",  x"0b",  x"a8",  x"f4",  x"93",  x"27",  x"8b", -- 1CE0
         x"00",  x"00",  x"1e",  x"01",  x"0b",  x"00",  x"ae",  x"80", -- 1CE8
         x"28",  x"08",  x"11",  x"22",  x"b2",  x"21",  x"01",  x"7e", -- 1CF0
         x"af",  x"e8",  x"c9",  x"80",  x"00",  x"40",  x"00",  x"00", -- 1CF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1D98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1DF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1E98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1ED8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1EF8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F00
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F08
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F10
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F18
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F20
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F28
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F30
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F38
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F40
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F48
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F50
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F58
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F60
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F68
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F70
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F78
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F80
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F88
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F90
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1F98
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FA8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FB8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FC8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FD8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FE8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 1FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 1FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;

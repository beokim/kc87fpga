library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity os is
    generic(
        AddrWidth   : integer := 9
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end os;

architecture rtl of os is
    type rom512x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom512x8 := (
         x"c3",  x"03",  x"f0",  x"31",  x"00",  x"02",  x"11",  x"00", -- 0000
         x"02",  x"21",  x"29",  x"f0",  x"01",  x"0c",  x"00",  x"ed", -- 0008
         x"b0",  x"3e",  x"02",  x"ed",  x"47",  x"ed",  x"5e",  x"3c", -- 0010
         x"d3",  x"8a",  x"3e",  x"cf",  x"d3",  x"8a",  x"af",  x"d3", -- 0018
         x"8a",  x"d3",  x"88",  x"cd",  x"35",  x"f0",  x"c3",  x"26", -- 0020
         x"f0",  x"d3",  x"f0",  x"00",  x"00",  x"9c",  x"f0",  x"fd", -- 0028
         x"f0",  x"85",  x"f0",  x"e9",  x"f0",  x"f3",  x"f5",  x"cd", -- 0030
         x"49",  x"f0",  x"f1",  x"f5",  x"cd",  x"67",  x"f0",  x"3e", -- 0038
         x"83",  x"d3",  x"93",  x"af",  x"d3",  x"90",  x"f1",  x"fb", -- 0040
         x"c9",  x"3e",  x"03",  x"d3",  x"80",  x"d3",  x"82",  x"d3", -- 0048
         x"8a",  x"af",  x"d3",  x"80",  x"3e",  x"c7",  x"d3",  x"83", -- 0050
         x"3e",  x"01",  x"d3",  x"83",  x"3e",  x"27",  x"d3",  x"82", -- 0058
         x"3e",  x"01",  x"d3",  x"82",  x"3e",  x"03",  x"c9",  x"3e", -- 0060
         x"cf",  x"d3",  x"92",  x"af",  x"d3",  x"92",  x"3e",  x"08", -- 0068
         x"d3",  x"93",  x"3e",  x"cf",  x"d3",  x"93",  x"3e",  x"ff", -- 0070
         x"d3",  x"93",  x"3e",  x"17",  x"d3",  x"93",  x"af",  x"d3", -- 0078
         x"93",  x"3d",  x"d3",  x"90",  x"c9",  x"f5",  x"3e",  x"0a", -- 0080
         x"32",  x"23",  x"00",  x"3e",  x"7f",  x"32",  x"24",  x"00", -- 0088
         x"3e",  x"a5",  x"d3",  x"82",  x"3e",  x"01",  x"d3",  x"82", -- 0090
         x"f1",  x"fb",  x"ed",  x"4d",  x"fb",  x"f5",  x"e5",  x"21", -- 0098
         x"23",  x"00",  x"35",  x"28",  x"13",  x"3e",  x"07",  x"a7", -- 00A0
         x"20",  x"21",  x"23",  x"cd",  x"d0",  x"f0",  x"28",  x"1b", -- 00A8
         x"bf",  x"28",  x"18",  x"2b",  x"36",  x"28",  x"18",  x"07", -- 00B0
         x"36",  x"06",  x"cd",  x"d0",  x"f0",  x"28",  x"0c",  x"23", -- 00B8
         x"77",  x"3a",  x"25",  x"00",  x"bf",  x"28",  x"04",  x"7e", -- 00C0
         x"32",  x"25",  x"00",  x"e1",  x"f1",  x"fb",  x"ed",  x"4d", -- 00C8
         x"3e",  x"20",  x"c9",  x"f5",  x"3e",  x"03",  x"d3",  x"80", -- 00D0
         x"3e",  x"85",  x"d3",  x"80",  x"3a",  x"6a",  x"00",  x"d3", -- 00D8
         x"80",  x"af",  x"32",  x"6a",  x"00",  x"f1",  x"fb",  x"ed", -- 00E0
         x"4d",  x"f5",  x"db",  x"80",  x"f5",  x"3e",  x"07",  x"d3", -- 00E8
         x"80",  x"3e",  x"b0",  x"d3",  x"80",  x"f1",  x"32",  x"6a", -- 00F0
         x"00",  x"f1",  x"fb",  x"ed",  x"4d",  x"fb",  x"e5",  x"c5", -- 00F8
         x"f5",  x"21",  x"20",  x"00",  x"06",  x"02",  x"3e",  x"3c", -- 0100
         x"2b",  x"34",  x"bf",  x"20",  x"0d",  x"36",  x"00",  x"10", -- 0108
         x"f7",  x"3e",  x"18",  x"2b",  x"34",  x"bf",  x"20",  x"02", -- 0110
         x"36",  x"00",  x"f1",  x"c1",  x"e1",  x"ed",  x"4d",  x"00", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0170
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0180
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0188
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0190
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0198
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 01F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity os is
    generic(
        AddrWidth   : integer := 12
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(AddrWidth-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end os;

architecture rtl of os is
    signal romAddr : integer range 0 to 2**AddrWidth-1;
    type rom4096x8 is array (0 to 2**AddrWidth-1) of std_logic_vector(7 downto 0); 
    constant romData : rom4096x8 := (
         x"c3",  x"64",  x"f6",  x"c3",  x"ae",  x"f6",  x"c3",  x"56", -- 0000
         x"f7",  x"c3",  x"7f",  x"f7",  x"c3",  x"83",  x"f7",  x"c3", -- 0008
         x"9e",  x"f7",  x"c3",  x"ae",  x"f7",  x"c3",  x"a8",  x"f7", -- 0010
         x"c3",  x"c4",  x"f7",  x"c3",  x"de",  x"f5",  x"c3",  x"0b", -- 0018
         x"f8",  x"c3",  x"fc",  x"f7",  x"c3",  x"df",  x"f7",  x"c3", -- 0020
         x"34",  x"f4",  x"c3",  x"6f",  x"f4",  x"c3",  x"a4",  x"f7", -- 0028
         x"c3",  x"33",  x"f7",  x"c3",  x"37",  x"f7",  x"c3",  x"de", -- 0030
         x"f5",  x"c3",  x"d2",  x"f7",  x"c3",  x"d9",  x"f7",  x"c3", -- 0038
         x"e5",  x"f7",  x"c3",  x"f4",  x"f7",  x"64",  x"f6",  x"09", -- 0040
         x"f0",  x"0c",  x"f0",  x"15",  x"f0",  x"12",  x"f0",  x"0f", -- 0048
         x"f0",  x"18",  x"f0",  x"39",  x"f0",  x"3c",  x"f0",  x"e2", -- 0050
         x"f3",  x"65",  x"f3",  x"06",  x"f0",  x"f3",  x"f3",  x"f8", -- 0058
         x"f3",  x"2d",  x"f4",  x"45",  x"f4",  x"6a",  x"f4",  x"3c", -- 0060
         x"f7",  x"3b",  x"f7",  x"de",  x"f5",  x"27",  x"f0",  x"2a", -- 0068
         x"f0",  x"1e",  x"f0",  x"21",  x"f0",  x"a8",  x"f4",  x"e3", -- 0070
         x"fa",  x"24",  x"f0",  x"3f",  x"f0",  x"42",  x"f0",  x"3e", -- 0078
         x"f7",  x"3d",  x"f7",  x"b9",  x"f5",  x"de",  x"f5",  x"d8", -- 0080
         x"f4",  x"21",  x"89",  x"f0",  x"e5",  x"21",  x"80",  x"00", -- 0088
         x"22",  x"1b",  x"00",  x"3e",  x"3e",  x"cd",  x"05",  x"f3", -- 0090
         x"cd",  x"5c",  x"f3",  x"38",  x"23",  x"cd",  x"b9",  x"f5", -- 0098
         x"d8",  x"21",  x"ea",  x"f5",  x"e5",  x"cd",  x"ea",  x"f1", -- 00A0
         x"ca",  x"e6",  x"f5",  x"c5",  x"cd",  x"8e",  x"f2",  x"c1", -- 00A8
         x"28",  x"07",  x"cd",  x"26",  x"f5",  x"d8",  x"2a",  x"71", -- 00B0
         x"00",  x"e9",  x"08",  x"30",  x"2a",  x"cd",  x"fe",  x"f2", -- 00B8
         x"da",  x"ae",  x"f6",  x"06",  x"04",  x"21",  x"e9",  x"ef", -- 00C0
         x"11",  x"d5",  x"fb",  x"cd",  x"e2",  x"f3",  x"3e",  x"3a", -- 00C8
         x"cd",  x"05",  x"f3",  x"d5",  x"5e",  x"23",  x"56",  x"23", -- 00D0
         x"e5",  x"cd",  x"e2",  x"f3",  x"e1",  x"d1",  x"13",  x"13", -- 00D8
         x"13",  x"cd",  x"fe",  x"f2",  x"10",  x"e5",  x"c9",  x"cd", -- 00E0
         x"ea",  x"f1",  x"28",  x"2c",  x"08",  x"da",  x"e6",  x"f5", -- 00E8
         x"c5",  x"01",  x"09",  x"04",  x"21",  x"d5",  x"fb",  x"cd", -- 00F0
         x"b8",  x"f2",  x"58",  x"c1",  x"20",  x"50",  x"3e",  x"04", -- 00F8
         x"93",  x"87",  x"32",  x"33",  x"00",  x"22",  x"40",  x"00", -- 0100
         x"79",  x"fe",  x"3a",  x"20",  x"05",  x"cd",  x"c4",  x"f1", -- 0108
         x"fe",  x"3d",  x"c2",  x"e2",  x"f5",  x"cd",  x"ea",  x"f1", -- 0110
         x"28",  x"5b",  x"c5",  x"cd",  x"b2",  x"f2",  x"c1",  x"28", -- 0118
         x"17",  x"cd",  x"ab",  x"f0",  x"d8",  x"00",  x"e5",  x"d5", -- 0120
         x"7c",  x"84",  x"85",  x"87",  x"16",  x"00",  x"5f",  x"21", -- 0128
         x"c9",  x"ef",  x"19",  x"71",  x"23",  x"70",  x"d1",  x"e1", -- 0130
         x"3a",  x"04",  x"00",  x"08",  x"30",  x"37",  x"3a",  x"33", -- 0138
         x"00",  x"47",  x"4d",  x"bc",  x"28",  x"0a",  x"95",  x"3c", -- 0140
         x"fe",  x"06",  x"28",  x"04",  x"3d",  x"b8",  x"20",  x"25", -- 0148
         x"d5",  x"58",  x"21",  x"04",  x"00",  x"06",  x"09",  x"3c", -- 0150
         x"cb",  x"1e",  x"3d",  x"20",  x"07",  x"cb",  x"39",  x"cb", -- 0158
         x"1e",  x"cb",  x"39",  x"05",  x"10",  x"f2",  x"43",  x"cd", -- 0160
         x"ce",  x"f2",  x"d1",  x"30",  x"0b",  x"08",  x"32",  x"04", -- 0168
         x"00",  x"3e",  x"04",  x"37",  x"c9",  x"c3",  x"e6",  x"f5", -- 0170
         x"2a",  x"40",  x"00",  x"73",  x"23",  x"72",  x"c3",  x"bd", -- 0178
         x"f0",  x"08",  x"38",  x"34",  x"06",  x"03",  x"3e",  x"17", -- 0180
         x"32",  x"2f",  x"00",  x"c5",  x"cd",  x"ea",  x"f1",  x"c1", -- 0188
         x"20",  x"e3",  x"d8",  x"5f",  x"3a",  x"2f",  x"00",  x"bb", -- 0190
         x"3e",  x"03",  x"d8",  x"4d",  x"6c",  x"63",  x"08",  x"38", -- 0198
         x"10",  x"3e",  x"3b",  x"10",  x"e3",  x"c3",  x"e2",  x"f5", -- 01A0
         x"22",  x"1e",  x"00",  x"79",  x"32",  x"1d",  x"00",  x"b7", -- 01A8
         x"c9",  x"1e",  x"00",  x"08",  x"10",  x"e5",  x"18",  x"f0", -- 01B0
         x"11",  x"01",  x"01",  x"cd",  x"a8",  x"f4",  x"cd",  x"e2", -- 01B8
         x"f3",  x"c3",  x"fe",  x"f2",  x"21",  x"81",  x"00",  x"23", -- 01C0
         x"7e",  x"fe",  x"20",  x"28",  x"fa",  x"cd",  x"d7",  x"f1", -- 01C8
         x"4f",  x"c0",  x"fe",  x"01",  x"d8",  x"bf",  x"c9",  x"7e", -- 01D0
         x"b7",  x"c8",  x"e5",  x"c5",  x"21",  x"ab",  x"fc",  x"01", -- 01D8
         x"05",  x"00",  x"ed",  x"b1",  x"c1",  x"e1",  x"36",  x"20", -- 01E0
         x"23",  x"c9",  x"11",  x"52",  x"01",  x"af",  x"06",  x"51", -- 01E8
         x"12",  x"1b",  x"10",  x"fc",  x"e5",  x"cd",  x"c4",  x"f1", -- 01F0
         x"38",  x"0d",  x"28",  x"0b",  x"12",  x"04",  x"13",  x"cd", -- 01F8
         x"d7",  x"f1",  x"20",  x"f8",  x"cd",  x"d0",  x"f1",  x"78", -- 0200
         x"32",  x"00",  x"01",  x"79",  x"e1",  x"08",  x"3a",  x"01", -- 0208
         x"01",  x"fe",  x"30",  x"38",  x"16",  x"fe",  x"3a",  x"30", -- 0210
         x"12",  x"e5",  x"c5",  x"11",  x"00",  x"01",  x"cd",  x"15", -- 0218
         x"f8",  x"c1",  x"e1",  x"38",  x"02",  x"bf",  x"c9",  x"bf", -- 0220
         x"c3",  x"e2",  x"f5",  x"fe",  x"40",  x"38",  x"f8",  x"37", -- 0228
         x"c9",  x"e5",  x"c5",  x"cd",  x"4d",  x"f2",  x"f5",  x"cb", -- 0230
         x"39",  x"18",  x"06",  x"e5",  x"c5",  x"cd",  x"4d",  x"f2", -- 0238
         x"f5",  x"cd",  x"69",  x"f2",  x"f1",  x"c1",  x"e1",  x"f5", -- 0240
         x"b7",  x"ed",  x"52",  x"f1",  x"c9",  x"11",  x"00",  x"04", -- 0248
         x"af",  x"ed",  x"52",  x"3c",  x"30",  x"fb",  x"21",  x"c1", -- 0250
         x"ef",  x"d6",  x"08",  x"23",  x"30",  x"fb",  x"c6",  x"08", -- 0258
         x"2b",  x"28",  x"fb",  x"06",  x"09",  x"cb",  x"16",  x"3d", -- 0260
         x"c8",  x"10",  x"fa",  x"c9",  x"e5",  x"d5",  x"eb",  x"1a", -- 0268
         x"fe",  x"20",  x"28",  x"04",  x"fe",  x"40",  x"38",  x"02", -- 0270
         x"e6",  x"df",  x"be",  x"13",  x"23",  x"20",  x"0c",  x"10", -- 0278
         x"ee",  x"d1",  x"d1",  x"6b",  x"62",  x"2b",  x"7e",  x"2b", -- 0280
         x"6e",  x"67",  x"c9",  x"d1",  x"e1",  x"c9",  x"21",  x"00", -- 0288
         x"fc",  x"e5",  x"3e",  x"c3",  x"ed",  x"a1",  x"20",  x"12", -- 0290
         x"23",  x"23",  x"c5",  x"01",  x"0b",  x"01",  x"cd",  x"b8", -- 0298
         x"f2",  x"c1",  x"28",  x"0c",  x"af",  x"2b",  x"2b",  x"be", -- 02A0
         x"20",  x"e8",  x"e1",  x"25",  x"20",  x"e3",  x"24",  x"c9", -- 02A8
         x"c1",  x"c9",  x"01",  x"06",  x"02",  x"21",  x"26",  x"fc", -- 02B0
         x"11",  x"01",  x"01",  x"c5",  x"41",  x"05",  x"05",  x"cd", -- 02B8
         x"6c",  x"f2",  x"c1",  x"c8",  x"79",  x"23",  x"3d",  x"20", -- 02C0
         x"fc",  x"10",  x"f0",  x"f6",  x"01",  x"c9",  x"f5",  x"16", -- 02C8
         x"00",  x"58",  x"78",  x"b7",  x"3a",  x"04",  x"00",  x"28", -- 02D0
         x"04",  x"cb",  x"3f",  x"10",  x"fc",  x"cb",  x"23",  x"e6", -- 02D8
         x"03",  x"83",  x"5f",  x"21",  x"c9",  x"ef",  x"f1",  x"19", -- 02E0
         x"19",  x"e5",  x"5e",  x"23",  x"56",  x"21",  x"ff",  x"ff", -- 02E8
         x"eb",  x"cd",  x"bc",  x"fc",  x"d1",  x"3f",  x"c9",  x"e5", -- 02F0
         x"d5",  x"c5",  x"ed",  x"b0",  x"18",  x"0e",  x"3e",  x"0d", -- 02F8
         x"cd",  x"05",  x"f3",  x"3e",  x"0a",  x"e5",  x"d5",  x"c5", -- 0300
         x"4f",  x"cd",  x"83",  x"f7",  x"c1",  x"d1",  x"e1",  x"c9", -- 0308
         x"3e",  x"20",  x"18",  x"f1",  x"ed",  x"73",  x"0b",  x"00", -- 0310
         x"31",  x"c0",  x"01",  x"37",  x"3f",  x"e5",  x"d5",  x"f5", -- 0318
         x"ed",  x"43",  x"0d",  x"00",  x"32",  x"0f",  x"00",  x"21", -- 0320
         x"45",  x"f3",  x"e5",  x"3e",  x"21",  x"b9",  x"da",  x"de", -- 0328
         x"f5",  x"06",  x"00",  x"21",  x"45",  x"f0",  x"09",  x"09", -- 0330
         x"7e",  x"23",  x"66",  x"6f",  x"4b",  x"42",  x"3a",  x"0f", -- 0338
         x"00",  x"e5",  x"2e",  x"03",  x"c9",  x"30",  x"06",  x"cd", -- 0340
         x"ea",  x"f5",  x"f1",  x"37",  x"f5",  x"f1",  x"d1",  x"e1", -- 0348
         x"3a",  x"0f",  x"00",  x"ed",  x"4b",  x"0d",  x"00",  x"ed", -- 0350
         x"7b",  x"0b",  x"00",  x"c9",  x"11",  x"80",  x"00",  x"3e", -- 0358
         x"50",  x"12",  x"3a",  x"0f",  x"00",  x"6b",  x"62",  x"23", -- 0360
         x"4d",  x"44",  x"03",  x"36",  x"00",  x"32",  x"35",  x"00", -- 0368
         x"e5",  x"d5",  x"c5",  x"cd",  x"7f",  x"f7",  x"c1",  x"d1", -- 0370
         x"e1",  x"d8",  x"e5",  x"21",  x"17",  x"00",  x"34",  x"35", -- 0378
         x"e1",  x"20",  x"2b",  x"fe",  x"03",  x"20",  x"03",  x"af", -- 0380
         x"37",  x"c9",  x"fe",  x"1f",  x"28",  x"1b",  x"fe",  x"02", -- 0388
         x"20",  x"07",  x"cd",  x"c6",  x"f3",  x"20",  x"fb",  x"18", -- 0390
         x"d7",  x"fe",  x"0d",  x"28",  x"20",  x"fe",  x"0b",  x"28", -- 0398
         x"cf",  x"fe",  x"0a",  x"28",  x"cb",  x"fe",  x"08",  x"20", -- 03A0
         x"05",  x"cd",  x"c6",  x"f3",  x"18",  x"c2",  x"fe",  x"10", -- 03A8
         x"28",  x"03",  x"34",  x"02",  x"03",  x"cd",  x"05",  x"f3", -- 03B0
         x"d8",  x"1a",  x"be",  x"20",  x"b3",  x"3a",  x"35",  x"00", -- 03B8
         x"32",  x"0f",  x"00",  x"c3",  x"fe",  x"f2",  x"34",  x"35", -- 03C0
         x"c8",  x"0b",  x"0a",  x"fe",  x"09",  x"28",  x"0c",  x"fe", -- 03C8
         x"20",  x"38",  x"f4",  x"3e",  x"08",  x"cd",  x"05",  x"f3", -- 03D0
         x"cd",  x"10",  x"f3",  x"3e",  x"08",  x"cd",  x"05",  x"f3", -- 03D8
         x"35",  x"c9",  x"1a",  x"b7",  x"20",  x"06",  x"3a",  x"17", -- 03E0
         x"00",  x"b7",  x"c8",  x"af",  x"cd",  x"05",  x"f3",  x"d8", -- 03E8
         x"13",  x"18",  x"ef",  x"21",  x"03",  x"01",  x"18",  x"38", -- 03F0
         x"cd",  x"93",  x"f5",  x"3c",  x"d8",  x"e5",  x"af",  x"32", -- 03F8
         x"6c",  x"00",  x"cd",  x"34",  x"f4",  x"e1",  x"22",  x"1b", -- 0400
         x"00",  x"d8",  x"e5",  x"11",  x"11",  x"00",  x"19",  x"11", -- 0408
         x"6d",  x"00",  x"01",  x"08",  x"00",  x"ed",  x"b0",  x"d1", -- 0410
         x"21",  x"5c",  x"00",  x"06",  x"0b",  x"cd",  x"6c",  x"f2", -- 0418
         x"3e",  x"0d",  x"37",  x"c0",  x"3a",  x"73",  x"00",  x"b7", -- 0420
         x"c8",  x"32",  x"c0",  x"ef",  x"c9",  x"21",  x"6d",  x"00", -- 0428
         x"22",  x"0d",  x"00",  x"c9",  x"cd",  x"d8",  x"f4",  x"d8", -- 0430
         x"22",  x"1b",  x"00",  x"21",  x"6c",  x"00",  x"34",  x"f5", -- 0438
         x"cd",  x"10",  x"f3",  x"f1",  x"c9",  x"cd",  x"93",  x"f5", -- 0440
         x"3c",  x"d8",  x"e5",  x"21",  x"5c",  x"00",  x"22",  x"1b", -- 0448
         x"00",  x"3e",  x"00",  x"32",  x"73",  x"00",  x"01",  x"70", -- 0450
         x"17",  x"af",  x"32",  x"6b",  x"00",  x"3e",  x"02",  x"32", -- 0458
         x"6c",  x"00",  x"cd",  x"72",  x"f4",  x"e1",  x"22",  x"1b", -- 0460
         x"00",  x"c9",  x"3e",  x"ff",  x"32",  x"6b",  x"00",  x"01", -- 0468
         x"a0",  x"00",  x"ed",  x"5b",  x"1b",  x"00",  x"3a",  x"c0", -- 0470
         x"ef",  x"b7",  x"28",  x"04",  x"3e",  x"09",  x"37",  x"c9", -- 0478
         x"2a",  x"36",  x"00",  x"d5",  x"11",  x"7f",  x"00",  x"ed", -- 0480
         x"52",  x"d1",  x"cd",  x"bc",  x"fc",  x"3e",  x"0a",  x"38", -- 0488
         x"ed",  x"eb",  x"cd",  x"3b",  x"f2",  x"30",  x"e5",  x"cd", -- 0490
         x"d6",  x"fe",  x"22",  x"1b",  x"00",  x"21",  x"6b",  x"00", -- 0498
         x"7e",  x"32",  x"0f",  x"00",  x"34",  x"c3",  x"e3",  x"fa", -- 04A0
         x"d5",  x"01",  x"1d",  x"00",  x"16",  x"03",  x"21",  x"01", -- 04A8
         x"01",  x"e5",  x"2b",  x"36",  x"3a",  x"23",  x"0a",  x"c5", -- 04B0
         x"b7",  x"28",  x"07",  x"47",  x"af",  x"c6",  x"01",  x"27", -- 04B8
         x"10",  x"fb",  x"77",  x"3e",  x"33",  x"ed",  x"67",  x"23", -- 04C0
         x"77",  x"23",  x"36",  x"00",  x"c1",  x"03",  x"15",  x"20", -- 04C8
         x"e2",  x"e1",  x"d1",  x"0e",  x"08",  x"c3",  x"f7",  x"f2", -- 04D0
         x"2a",  x"36",  x"00",  x"11",  x"7f",  x"00",  x"ed",  x"52", -- 04D8
         x"ed",  x"5b",  x"1b",  x"00",  x"cd",  x"bc",  x"fc",  x"3e", -- 04E0
         x"0a",  x"d8",  x"eb",  x"cd",  x"3b",  x"f2",  x"3e",  x"09", -- 04E8
         x"30",  x"1d",  x"f5",  x"f1",  x"cd",  x"59",  x"ff",  x"cd", -- 04F0
         x"e3",  x"fa",  x"f5",  x"e5",  x"21",  x"6c",  x"00",  x"3a", -- 04F8
         x"6b",  x"00",  x"be",  x"e1",  x"38",  x"ed",  x"28",  x"09", -- 0500
         x"fe",  x"ff",  x"28",  x"05",  x"f1",  x"3e",  x"0b",  x"37", -- 0508
         x"c9",  x"f1",  x"3e",  x"0c",  x"d8",  x"3a",  x"6b",  x"00", -- 0510
         x"3c",  x"3e",  x"00",  x"20",  x"01",  x"3c",  x"32",  x"0f", -- 0518
         x"00",  x"c9",  x"cd",  x"ea",  x"f1",  x"c8",  x"21",  x"e6", -- 0520
         x"f5",  x"e5",  x"3a",  x"00",  x"01",  x"fe",  x"09",  x"d0", -- 0528
         x"11",  x"5c",  x"00",  x"3e",  x"08",  x"cd",  x"88",  x"f5", -- 0530
         x"08",  x"30",  x"0e",  x"08",  x"21",  x"43",  x"4f",  x"22", -- 0538
         x"64",  x"00",  x"3e",  x"4d",  x"32",  x"66",  x"00",  x"18", -- 0540
         x"16",  x"79",  x"fe",  x"2e",  x"e1",  x"c2",  x"e2",  x"f5", -- 0548
         x"e5",  x"cd",  x"ea",  x"f1",  x"c8",  x"3e",  x"03",  x"b8", -- 0550
         x"d8",  x"11",  x"64",  x"00",  x"cd",  x"88",  x"f5",  x"e1", -- 0558
         x"08",  x"d2",  x"e2",  x"f5",  x"cd",  x"f8",  x"f3",  x"30", -- 0560
         x"09",  x"b7",  x"37",  x"c8",  x"cd",  x"a3",  x"f5",  x"d8", -- 0568
         x"18",  x"f2",  x"2a",  x"6d",  x"00",  x"22",  x"1b",  x"00", -- 0570
         x"cd",  x"34",  x"f4",  x"30",  x"05",  x"cd",  x"a3",  x"f5", -- 0578
         x"d8",  x"af",  x"b7",  x"28",  x"f3",  x"c3",  x"fe",  x"f2", -- 0580
         x"21",  x"01",  x"01",  x"47",  x"7e",  x"12",  x"23",  x"13", -- 0588
         x"10",  x"fa",  x"c9",  x"11",  x"48",  x"fc",  x"cd",  x"e2", -- 0590
         x"f3",  x"cd",  x"5c",  x"f3",  x"2a",  x"1b",  x"00",  x"d0", -- 0598
         x"3e",  x"ff",  x"c9",  x"cd",  x"ea",  x"f5",  x"cd",  x"99", -- 05A0
         x"f5",  x"d8",  x"3a",  x"0f",  x"00",  x"fe",  x"09",  x"37", -- 05A8
         x"3f",  x"c0",  x"0e",  x"01",  x"cd",  x"31",  x"f2",  x"b7", -- 05B0
         x"c9",  x"13",  x"1a",  x"b7",  x"28",  x"1e",  x"6b",  x"62", -- 05B8
         x"e5",  x"23",  x"13",  x"47",  x"0e",  x"00",  x"eb",  x"3e", -- 05C0
         x"1f",  x"be",  x"30",  x"05",  x"ed",  x"a0",  x"03",  x"03", -- 05C8
         x"2b",  x"23",  x"10",  x"f5",  x"e1",  x"71",  x"eb",  x"79", -- 05D0
         x"b7",  x"36",  x"00",  x"c0",  x"37",  x"c9",  x"3e",  x"07", -- 05D8
         x"37",  x"c9",  x"3e",  x"02",  x"37",  x"c9",  x"3e",  x"01", -- 05E0
         x"37",  x"c9",  x"d0",  x"fe",  x"ff",  x"37",  x"c8",  x"32", -- 05E8
         x"0f",  x"00",  x"b7",  x"37",  x"c8",  x"f5",  x"af",  x"32", -- 05F0
         x"15",  x"00",  x"cd",  x"fe",  x"f2",  x"f1",  x"11",  x"5b", -- 05F8
         x"fc",  x"d6",  x"05",  x"30",  x"0c",  x"f5",  x"cd",  x"e2", -- 0600
         x"f3",  x"f1",  x"c6",  x"35",  x"cd",  x"05",  x"f3",  x"18", -- 0608
         x"4d",  x"d6",  x"02",  x"d8",  x"f5",  x"11",  x"56",  x"fc", -- 0610
         x"cd",  x"e2",  x"f3",  x"3e",  x"3a",  x"cd",  x"05",  x"f3", -- 0618
         x"cd",  x"10",  x"f3",  x"f1",  x"20",  x"04",  x"06",  x"08", -- 0620
         x"18",  x"03",  x"3d",  x"20",  x"0f",  x"21",  x"cc",  x"fb", -- 0628
         x"11",  x"09",  x"00",  x"cb",  x"38",  x"04",  x"19",  x"10", -- 0630
         x"fd",  x"eb",  x"18",  x"1f",  x"11",  x"62",  x"fc",  x"3d", -- 0638
         x"28",  x"19",  x"11",  x"73",  x"fc",  x"3d",  x"28",  x"13", -- 0640
         x"11",  x"81",  x"fc",  x"3d",  x"28",  x"0d",  x"11",  x"92", -- 0648
         x"fc",  x"3d",  x"28",  x"07",  x"11",  x"9d",  x"fc",  x"3d", -- 0650
         x"28",  x"01",  x"1b",  x"cd",  x"e2",  x"f3",  x"cd",  x"fe", -- 0658
         x"f2",  x"af",  x"37",  x"c9",  x"f3",  x"31",  x"00",  x"02", -- 0660
         x"0e",  x"00",  x"2a",  x"36",  x"00",  x"5d",  x"54",  x"13", -- 0668
         x"06",  x"01",  x"ed",  x"b0",  x"3e",  x"02",  x"ed",  x"47", -- 0670
         x"3c",  x"d3",  x"8a",  x"3e",  x"cf",  x"d3",  x"8a",  x"af", -- 0678
         x"d3",  x"8a",  x"d3",  x"88",  x"21",  x"c1",  x"ef",  x"3e", -- 0680
         x"ff",  x"77",  x"23",  x"77",  x"23",  x"3c",  x"06",  x"05", -- 0688
         x"77",  x"23",  x"10",  x"fc",  x"3e",  x"30",  x"77",  x"00", -- 0690
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"21", -- 0698
         x"14",  x"f3",  x"22",  x"06",  x"00",  x"cd",  x"e0",  x"f6", -- 06A0
         x"11",  x"30",  x"fc",  x"cd",  x"e2",  x"f3",  x"f3",  x"31", -- 06A8
         x"00",  x"02",  x"3e",  x"c3",  x"32",  x"00",  x"00",  x"32", -- 06B0
         x"05",  x"00",  x"21",  x"ae",  x"f6",  x"22",  x"01",  x"00", -- 06B8
         x"3a",  x"04",  x"00",  x"e6",  x"fc",  x"f6",  x"01",  x"cd", -- 06C0
         x"12",  x"f7",  x"11",  x"f7",  x"fb",  x"cd",  x"e2",  x"f3", -- 06C8
         x"21",  x"23",  x"00",  x"22",  x"82",  x"00",  x"cd",  x"ea", -- 06D0
         x"f1",  x"cd",  x"8e",  x"f2",  x"c2",  x"89",  x"f0",  x"e9", -- 06D8
         x"21",  x"c9",  x"ef",  x"11",  x"ca",  x"ef",  x"01",  x"1f", -- 06E0
         x"00",  x"36",  x"ff",  x"ed",  x"b0",  x"11",  x"00",  x"02", -- 06E8
         x"21",  x"b0",  x"fc",  x"0e",  x"0c",  x"ed",  x"b0",  x"21", -- 06F0
         x"24",  x"fc",  x"22",  x"eb",  x"ef",  x"22",  x"ed",  x"ef", -- 06F8
         x"22",  x"ef",  x"ef",  x"21",  x"b4",  x"f7",  x"22",  x"cd", -- 0700
         x"ef",  x"af",  x"32",  x"27",  x"00",  x"32",  x"c0",  x"ef", -- 0708
         x"3e",  x"01",  x"32",  x"04",  x"00",  x"21",  x"26",  x"fc", -- 0710
         x"22",  x"e9",  x"ef",  x"21",  x"f1",  x"f8",  x"22",  x"cb", -- 0718
         x"ef",  x"22",  x"e3",  x"ef",  x"ed",  x"5e",  x"11",  x"ff", -- 0720
         x"ff",  x"1b",  x"7b",  x"b2",  x"00",  x"00",  x"32",  x"15", -- 0728
         x"00",  x"3d",  x"e9",  x"2e",  x"07",  x"18",  x"07",  x"2e", -- 0730
         x"05",  x"59",  x"50",  x"2c",  x"2c",  x"2c",  x"7d",  x"cd", -- 0738
         x"58",  x"f7",  x"d8",  x"fe",  x"03",  x"c8",  x"4d",  x"44", -- 0740
         x"fe",  x"06",  x"d0",  x"22",  x"0d",  x"00",  x"fe",  x"04", -- 0748
         x"c8",  x"ed",  x"53",  x"bc",  x"01",  x"c9",  x"3e",  x"00", -- 0750
         x"06",  x"00",  x"c5",  x"d5",  x"cd",  x"ce",  x"f2",  x"d1", -- 0758
         x"30",  x"04",  x"c1",  x"3e",  x"08",  x"c9",  x"e5",  x"21", -- 0760
         x"6f",  x"f7",  x"e3",  x"32",  x"2f",  x"00",  x"e9",  x"c1", -- 0768
         x"4f",  x"38",  x"f0",  x"3a",  x"2f",  x"00",  x"fe",  x"02", -- 0770
         x"d0",  x"79",  x"32",  x"0f",  x"00",  x"b7",  x"c9",  x"3e", -- 0778
         x"01",  x"18",  x"d5",  x"79",  x"fe",  x"10",  x"20",  x"08", -- 0780
         x"3a",  x"15",  x"00",  x"ee",  x"01",  x"32",  x"15",  x"00", -- 0788
         x"3e",  x"02",  x"c5",  x"cd",  x"58",  x"f7",  x"e1",  x"4d", -- 0790
         x"d8",  x"3a",  x"15",  x"00",  x"b7",  x"c8",  x"3e",  x"02", -- 0798
         x"06",  x"06",  x"18",  x"b6",  x"3e",  x"00",  x"18",  x"f8", -- 07A0
         x"3e",  x"01",  x"06",  x"02",  x"18",  x"ac",  x"3e",  x"02", -- 07A8
         x"06",  x"04",  x"18",  x"a6",  x"fe",  x"01",  x"28",  x"f0", -- 07B0
         x"fe",  x"ff",  x"20",  x"e4",  x"cd",  x"aa",  x"f7",  x"d8", -- 07B8
         x"3e",  x"ff",  x"18",  x"dc",  x"cd",  x"8f",  x"fe",  x"ed", -- 07C0
         x"4b",  x"13",  x"00",  x"ed",  x"43",  x"0d",  x"00",  x"c3", -- 07C8
         x"e9",  x"fa",  x"3a",  x"04",  x"00",  x"32",  x"0f",  x"00", -- 07D0
         x"4f",  x"79",  x"32",  x"04",  x"00",  x"b7",  x"c9",  x"ed", -- 07D8
         x"43",  x"1b",  x"00",  x"b7",  x"c9",  x"69",  x"60",  x"cd", -- 07E0
         x"3b",  x"f2",  x"3e",  x"01",  x"38",  x"01",  x"3d",  x"32", -- 07E8
         x"0f",  x"00",  x"b7",  x"c9",  x"69",  x"60",  x"4f",  x"cd", -- 07F0
         x"31",  x"f2",  x"b7",  x"c9",  x"3a",  x"1d",  x"00",  x"32", -- 07F8
         x"0f",  x"00",  x"2a",  x"1e",  x"00",  x"4c",  x"45",  x"ed", -- 0800
         x"43",  x"0d",  x"00",  x"32",  x"1d",  x"00",  x"68",  x"61", -- 0808
         x"22",  x"1e",  x"00",  x"b7",  x"c9",  x"1a",  x"b7",  x"37", -- 0810
         x"c8",  x"3e",  x"02",  x"cd",  x"36",  x"f8",  x"d8",  x"01", -- 0818
         x"02",  x"00",  x"1a",  x"13",  x"d6",  x"30",  x"d8",  x"fe", -- 0820
         x"0a",  x"3f",  x"d8",  x"80",  x"0d",  x"c8",  x"87",  x"47", -- 0828
         x"87",  x"87",  x"80",  x"47",  x"18",  x"ec",  x"6b",  x"62", -- 0830
         x"13",  x"be",  x"c8",  x"06",  x"00",  x"4e",  x"38",  x"13", -- 0838
         x"77",  x"91",  x"09",  x"5d",  x"54",  x"13",  x"c5",  x"ed", -- 0840
         x"b8",  x"c1",  x"eb",  x"36",  x"30",  x"eb",  x"03",  x"3d", -- 0848
         x"20",  x"f0",  x"c9",  x"f5",  x"23",  x"23",  x"1a",  x"fe", -- 0850
         x"30",  x"20",  x"0a",  x"0d",  x"cd",  x"f7",  x"f2",  x"1b", -- 0858
         x"79",  x"12",  x"f1",  x"18",  x"d1",  x"f1",  x"37",  x"c9", -- 0860
         x"d6",  x"14",  x"38",  x"15",  x"28",  x"06",  x"06",  x"f8", -- 0868
         x"7b",  x"a0",  x"b1",  x"c9",  x"7b",  x"06",  x"8f",  x"cb", -- 0870
         x"21",  x"cb",  x"21",  x"cb",  x"21",  x"cb",  x"21",  x"18", -- 0878
         x"f0",  x"db",  x"88",  x"06",  x"c7",  x"cd",  x"79",  x"f8", -- 0880
         x"d3",  x"88",  x"f1",  x"18",  x"0e",  x"3a",  x"27",  x"00", -- 0888
         x"5f",  x"7e",  x"b7",  x"28",  x"09",  x"cd",  x"68",  x"f8", -- 0890
         x"32",  x"27",  x"00",  x"af",  x"77",  x"c9",  x"79",  x"d6", -- 0898
         x"05",  x"28",  x"39",  x"3d",  x"20",  x"05",  x"7b",  x"ee", -- 08A0
         x"80",  x"18",  x"ed",  x"3d",  x"20",  x"1d",  x"f3",  x"cd", -- 08A8
         x"c4",  x"f8",  x"cd",  x"0d",  x"ff",  x"01",  x"30",  x"00", -- 08B0
         x"cd",  x"31",  x"ff",  x"ed",  x"a1",  x"ea",  x"b8",  x"f8", -- 08B8
         x"3e",  x"03",  x"d3",  x"80",  x"db",  x"88",  x"ee",  x"80", -- 08C0
         x"d3",  x"88",  x"c9",  x"d6",  x"0a",  x"20",  x"06",  x"2b", -- 08C8
         x"7e",  x"ee",  x"01",  x"77",  x"c9",  x"d6",  x"03",  x"28", -- 08D0
         x"03",  x"3d",  x"20",  x"02",  x"79",  x"77",  x"3d",  x"28", -- 08D8
         x"0a",  x"cd",  x"7d",  x"f9",  x"3a",  x"16",  x"00",  x"b7", -- 08E0
         x"c8",  x"18",  x"c3",  x"7b",  x"cd",  x"d6",  x"fa",  x"18", -- 08E8
         x"a7",  x"21",  x"17",  x"00",  x"3c",  x"20",  x"23",  x"f3", -- 08F0
         x"21",  x"00",  x"19",  x"22",  x"3b",  x"00",  x"26",  x"29", -- 08F8
         x"22",  x"3d",  x"00",  x"26",  x"00",  x"22",  x"23",  x"00", -- 0900
         x"22",  x"25",  x"00",  x"22",  x"13",  x"00",  x"22",  x"16", -- 0908
         x"00",  x"db",  x"88",  x"e6",  x"38",  x"d3",  x"88",  x"c3", -- 0910
         x"e3",  x"fa",  x"3d",  x"20",  x"04",  x"3a",  x"25",  x"00", -- 0918
         x"c9",  x"3d",  x"20",  x"21",  x"3a",  x"25",  x"00",  x"b7", -- 0920
         x"28",  x"fa",  x"f5",  x"af",  x"32",  x"25",  x"00",  x"32", -- 0928
         x"13",  x"00",  x"32",  x"14",  x"00",  x"7e",  x"b7",  x"28", -- 0930
         x"0a",  x"f1",  x"fe",  x"39",  x"30",  x"e6",  x"d6",  x"31", -- 0938
         x"38",  x"e2",  x"f5",  x"f1",  x"c9",  x"3d",  x"ca",  x"8d", -- 0940
         x"f8",  x"0e",  x"00",  x"3d",  x"ca",  x"33",  x"fa",  x"3d", -- 0948
         x"ca",  x"f3",  x"f9",  x"3d",  x"20",  x"08",  x"cd",  x"7d", -- 0950
         x"f9",  x"ed",  x"5b",  x"2b",  x"00",  x"c9",  x"3d",  x"28", -- 0958
         x"18",  x"3d",  x"28",  x"19",  x"3d",  x"c0",  x"21",  x"00", -- 0960
         x"ec",  x"eb",  x"ed",  x"52",  x"d8",  x"11",  x"28",  x"00", -- 0968
         x"ed",  x"52",  x"3c",  x"30",  x"fb",  x"19",  x"2c",  x"67", -- 0970
         x"eb",  x"ed",  x"53",  x"2b",  x"00",  x"21",  x"f3",  x"f9", -- 0978
         x"e5",  x"cd",  x"33",  x"fa",  x"79",  x"d6",  x"08",  x"d8", -- 0980
         x"28",  x"4e",  x"3d",  x"28",  x"30",  x"3d",  x"28",  x"3b", -- 0988
         x"3d",  x"28",  x"53",  x"3d",  x"28",  x"0d",  x"3d",  x"28", -- 0990
         x"1e",  x"fe",  x"13",  x"d8",  x"71",  x"3a",  x"27",  x"00", -- 0998
         x"12",  x"18",  x"1a",  x"3a",  x"3b",  x"00",  x"3c",  x"32", -- 09A0
         x"2c",  x"00",  x"47",  x"3a",  x"3c",  x"00",  x"90",  x"47", -- 09A8
         x"c5",  x"cd",  x"4f",  x"fa",  x"c1",  x"10",  x"f9",  x"3a", -- 09B0
         x"3d",  x"00",  x"32",  x"2b",  x"00",  x"21",  x"2b",  x"00", -- 09B8
         x"11",  x"3e",  x"00",  x"34",  x"1a",  x"be",  x"c0",  x"1b", -- 09C0
         x"1a",  x"3c",  x"77",  x"21",  x"2c",  x"00",  x"34",  x"3a", -- 09C8
         x"3c",  x"00",  x"3d",  x"be",  x"d0",  x"77",  x"18",  x"77", -- 09D0
         x"21",  x"2b",  x"00",  x"11",  x"3d",  x"00",  x"35",  x"1a", -- 09D8
         x"be",  x"c0",  x"13",  x"1a",  x"3d",  x"77",  x"21",  x"2c", -- 09E0
         x"00",  x"35",  x"3a",  x"3b",  x"00",  x"be",  x"d8",  x"3c", -- 09E8
         x"77",  x"18",  x"5d",  x"3a",  x"2b",  x"00",  x"4f",  x"3a", -- 09F0
         x"2c",  x"00",  x"47",  x"21",  x"d8",  x"eb",  x"11",  x"28", -- 09F8
         x"00",  x"19",  x"10",  x"fd",  x"41",  x"2b",  x"23",  x"10", -- 0A00
         x"fd",  x"22",  x"2d",  x"00",  x"3a",  x"c8",  x"ef",  x"cb", -- 0A08
         x"6f",  x"20",  x"06",  x"7e",  x"32",  x"3f",  x"00",  x"36", -- 0A10
         x"ff",  x"11",  x"00",  x"04",  x"e5",  x"ed",  x"52",  x"7e", -- 0A18
         x"32",  x"34",  x"00",  x"3a",  x"27",  x"00",  x"ee",  x"80", -- 0A20
         x"47",  x"ae",  x"e6",  x"f0",  x"78",  x"cc",  x"d6",  x"fa", -- 0A28
         x"77",  x"e1",  x"c9",  x"2a",  x"2d",  x"00",  x"3a",  x"c8", -- 0A30
         x"ef",  x"cb",  x"6f",  x"20",  x"04",  x"3a",  x"3f",  x"00", -- 0A38
         x"77",  x"11",  x"00",  x"04",  x"e5",  x"b7",  x"ed",  x"52", -- 0A40
         x"3a",  x"34",  x"00",  x"77",  x"eb",  x"e1",  x"c9",  x"3e", -- 0A48
         x"af",  x"f5",  x"21",  x"d8",  x"eb",  x"11",  x"28",  x"00", -- 0A50
         x"3a",  x"3b",  x"00",  x"3c",  x"4f",  x"3a",  x"3c",  x"00", -- 0A58
         x"3d",  x"47",  x"f1",  x"c5",  x"b7",  x"28",  x"01",  x"41", -- 0A60
         x"19",  x"10",  x"fd",  x"c1",  x"f5",  x"78",  x"91",  x"28", -- 0A68
         x"37",  x"47",  x"f1",  x"e5",  x"b7",  x"28",  x"03",  x"19", -- 0A70
         x"18",  x"02",  x"ed",  x"52",  x"d1",  x"f5",  x"e5",  x"c5", -- 0A78
         x"3a",  x"3d",  x"00",  x"3c",  x"47",  x"2b",  x"1b",  x"23", -- 0A80
         x"13",  x"10",  x"fc",  x"4f",  x"3a",  x"3e",  x"00",  x"91", -- 0A88
         x"4f",  x"cd",  x"f7",  x"f2",  x"c5",  x"01",  x"00",  x"04", -- 0A90
         x"eb",  x"ed",  x"42",  x"eb",  x"ed",  x"42",  x"c1",  x"ed", -- 0A98
         x"b0",  x"c1",  x"e1",  x"11",  x"28",  x"00",  x"10",  x"ca", -- 0AA0
         x"f1",  x"3a",  x"3d",  x"00",  x"3c",  x"4f",  x"47",  x"23", -- 0AA8
         x"10",  x"fd",  x"5d",  x"54",  x"2b",  x"3a",  x"3e",  x"00", -- 0AB0
         x"91",  x"4f",  x"0d",  x"36",  x"20",  x"c5",  x"f5",  x"c4", -- 0AB8
         x"f7",  x"f2",  x"11",  x"00",  x"04",  x"ed",  x"52",  x"3a", -- 0AC0
         x"27",  x"00",  x"cb",  x"bf",  x"77",  x"f1",  x"c1",  x"c8", -- 0AC8
         x"5d",  x"54",  x"13",  x"ed",  x"b0",  x"c9",  x"0e",  x"00", -- 0AD0
         x"cb",  x"27",  x"cb",  x"19",  x"07",  x"07",  x"07",  x"e6", -- 0AD8
         x"7f",  x"b1",  x"c9",  x"f3",  x"f5",  x"cd",  x"f7",  x"fa", -- 0AE0
         x"f1",  x"f5",  x"cd",  x"15",  x"fb",  x"3e",  x"83",  x"d3", -- 0AE8
         x"93",  x"af",  x"d3",  x"90",  x"f1",  x"fb",  x"c9",  x"3e", -- 0AF0
         x"03",  x"d3",  x"80",  x"d3",  x"82",  x"d3",  x"8a",  x"af", -- 0AF8
         x"d3",  x"80",  x"3e",  x"c7",  x"d3",  x"83",  x"3e",  x"40", -- 0B00
         x"d3",  x"83",  x"3e",  x"27",  x"d3",  x"82",  x"3e",  x"96", -- 0B08
         x"d3",  x"82",  x"3e",  x"03",  x"c9",  x"3e",  x"cf",  x"d3", -- 0B10
         x"92",  x"af",  x"d3",  x"92",  x"3e",  x"08",  x"d3",  x"93", -- 0B18
         x"3e",  x"cf",  x"d3",  x"93",  x"3e",  x"ff",  x"d3",  x"93", -- 0B20
         x"3e",  x"17",  x"d3",  x"93",  x"af",  x"d3",  x"93",  x"3d", -- 0B28
         x"d3",  x"90",  x"c9",  x"18",  x"1e",  x"1f",  x"5d",  x"00", -- 0B30
         x"08",  x"09",  x"0a",  x"0b",  x"02",  x"0d",  x"03",  x"20", -- 0B38
         x"19",  x"13",  x"1a",  x"5e",  x"00",  x"08",  x"09",  x"0a", -- 0B40
         x"0b",  x"1b",  x"0d",  x"03",  x"20",  x"00",  x"14",  x"00", -- 0B48
         x"7e",  x"1c",  x"1d",  x"7d",  x"ab",  x"8d",  x"82",  x"85", -- 0B50
         x"86",  x"84",  x"cf",  x"c3",  x"96",  x"90",  x"9b",  x"9c", -- 0B58
         x"af",  x"c4",  x"95",  x"92",  x"ae",  x"87",  x"ac",  x"8c", -- 0B60
         x"91",  x"83",  x"ad",  x"80",  x"81",  x"c2",  x"00",  x"00", -- 0B68
         x"00",  x"93",  x"00",  x"00",  x"ec",  x"ed",  x"ee",  x"ef", -- 0B70
         x"f0",  x"ca",  x"cc",  x"d0",  x"d1",  x"da",  x"de",  x"fc", -- 0B78
         x"df",  x"fd",  x"db",  x"b3",  x"a0",  x"a1",  x"9e",  x"9f", -- 0B80
         x"c0",  x"c7",  x"b4",  x"b0",  x"b1",  x"8f",  x"fe",  x"dc", -- 0B88
         x"ff",  x"dd",  x"be",  x"b2",  x"a3",  x"f9",  x"aa",  x"a5", -- 0B90
         x"a9",  x"88",  x"c8",  x"c6",  x"bc",  x"b6",  x"bb",  x"ba", -- 0B98
         x"fb",  x"fa",  x"bd",  x"b8",  x"a8",  x"c1",  x"a6",  x"89", -- 0BA0
         x"b5",  x"f8",  x"a4",  x"a2",  x"a7",  x"c5",  x"98",  x"00", -- 0BA8
         x"d7",  x"b9",  x"d2",  x"d3",  x"f2",  x"e0",  x"e2",  x"f4", -- 0BB0
         x"e8",  x"f5",  x"f6",  x"8a",  x"d4",  x"8b",  x"d8",  x"d9", -- 0BB8
         x"cd",  x"ce",  x"d5",  x"d6",  x"ea",  x"e7",  x"f3",  x"e6", -- 0BC0
         x"c9",  x"e1",  x"e9",  x"e3",  x"e4",  x"cb",  x"94",  x"9d", -- 0BC8
         x"97",  x"9a",  x"99",  x"e9",  x"ef",  x"43",  x"4f",  x"4e", -- 0BD0
         x"53",  x"54",  x"20",  x"00",  x"eb",  x"ef",  x"52",  x"45", -- 0BD8
         x"41",  x"44",  x"45",  x"52",  x"00",  x"ed",  x"ef",  x"50", -- 0BE0
         x"55",  x"4e",  x"43",  x"48",  x"20",  x"00",  x"ef",  x"ef", -- 0BE8
         x"4c",  x"49",  x"53",  x"54",  x"20",  x"20",  x"00",  x"0a", -- 0BF0
         x"0d",  x"4f",  x"53",  x"0a",  x"0d",  x"00",  x"ff",  x"ff", -- 0BF8
         x"c3",  x"ba",  x"f0",  x"41",  x"53",  x"47",  x"4e",  x"20", -- 0C00
         x"20",  x"20",  x"20",  x"00",  x"c3",  x"81",  x"f1",  x"54", -- 0C08
         x"49",  x"4d",  x"45",  x"20",  x"20",  x"20",  x"20",  x"00", -- 0C10
         x"c3",  x"22",  x"f5",  x"43",  x"4c",  x"4f",  x"41",  x"44", -- 0C18
         x"20",  x"20",  x"20",  x"00",  x"01",  x"00",  x"43",  x"52", -- 0C20
         x"54",  x"00",  x"02",  x"00",  x"42",  x"41",  x"54",  x"00", -- 0C28
         x"14",  x"01",  x"0c",  x"72",  x"6f",  x"62",  x"6f",  x"74", -- 0C30
         x"72",  x"6f",  x"6e",  x"20",  x"20",  x"5a",  x"20",  x"39", -- 0C38
         x"30",  x"30",  x"31",  x"0a",  x"0d",  x"14",  x"02",  x"00", -- 0C40
         x"0a",  x"73",  x"74",  x"61",  x"72",  x"74",  x"20",  x"74", -- 0C48
         x"61",  x"70",  x"65",  x"0a",  x"0d",  x"00",  x"07",  x"42", -- 0C50
         x"4f",  x"53",  x"2d",  x"65",  x"72",  x"72",  x"6f",  x"72", -- 0C58
         x"07",  x"00",  x"6d",  x"65",  x"6d",  x"6f",  x"72",  x"79", -- 0C60
         x"20",  x"70",  x"72",  x"6f",  x"74",  x"65",  x"63",  x"74", -- 0C68
         x"65",  x"64",  x"00",  x"65",  x"6e",  x"64",  x"20",  x"6f", -- 0C70
         x"66",  x"20",  x"6d",  x"65",  x"6d",  x"6f",  x"72",  x"79", -- 0C78
         x"00",  x"72",  x"65",  x"63",  x"6f",  x"72",  x"64",  x"20", -- 0C80
         x"6e",  x"6f",  x"74",  x"20",  x"66",  x"6f",  x"75",  x"6e", -- 0C88
         x"64",  x"00",  x"62",  x"61",  x"64",  x"20",  x"72",  x"65", -- 0C90
         x"63",  x"6f",  x"72",  x"64",  x"00",  x"66",  x"69",  x"6c", -- 0C98
         x"65",  x"20",  x"6e",  x"6f",  x"74",  x"20",  x"66",  x"6f", -- 0CA0
         x"75",  x"6e",  x"64",  x"00",  x"20",  x"2c",  x"2e",  x"3a", -- 0CA8
         x"43",  x"ff",  x"00",  x"00",  x"fb",  x"fc",  x"c2",  x"fc", -- 0CB0
         x"e4",  x"fc",  x"bd",  x"ff",  x"e5",  x"b7",  x"ed",  x"52", -- 0CB8
         x"e1",  x"c9",  x"fb",  x"e5",  x"c5",  x"f5",  x"21",  x"20", -- 0CC0
         x"00",  x"06",  x"02",  x"3e",  x"3c",  x"2b",  x"34",  x"be", -- 0CC8
         x"20",  x"0d",  x"36",  x"00",  x"10",  x"f7",  x"3e",  x"18", -- 0CD0
         x"2b",  x"34",  x"be",  x"20",  x"02",  x"36",  x"00",  x"f1", -- 0CD8
         x"c1",  x"e1",  x"ed",  x"4d",  x"f5",  x"3e",  x"0a",  x"32", -- 0CE0
         x"23",  x"00",  x"3e",  x"7f",  x"32",  x"24",  x"00",  x"3e", -- 0CE8
         x"a5",  x"d3",  x"82",  x"3e",  x"01",  x"d3",  x"82",  x"f1", -- 0CF0
         x"fb",  x"ed",  x"4d",  x"fb",  x"f5",  x"e5",  x"21",  x"23", -- 0CF8
         x"00",  x"35",  x"28",  x"13",  x"3e",  x"07",  x"a6",  x"20", -- 0D00
         x"22",  x"23",  x"cd",  x"30",  x"fd",  x"28",  x"1c",  x"be", -- 0D08
         x"28",  x"19",  x"2b",  x"36",  x"28",  x"18",  x"07",  x"36", -- 0D10
         x"06",  x"cd",  x"33",  x"fd",  x"28",  x"0d",  x"23",  x"77", -- 0D18
         x"3a",  x"25",  x"00",  x"fe",  x"03",  x"28",  x"04",  x"7e", -- 0D20
         x"32",  x"25",  x"00",  x"e1",  x"f1",  x"fb",  x"ed",  x"4d", -- 0D28
         x"7e",  x"b7",  x"c8",  x"e5",  x"d5",  x"c5",  x"21",  x"68", -- 0D30
         x"fe",  x"e5",  x"cd",  x"8f",  x"fe",  x"7a",  x"b7",  x"c8", -- 0D38
         x"7b",  x"b7",  x"c8",  x"3a",  x"26",  x"00",  x"b7",  x"28", -- 0D40
         x"06",  x"cb",  x"c3",  x"cb",  x"fa",  x"cb",  x"bd",  x"e5", -- 0D48
         x"d5",  x"5a",  x"0e",  x"08",  x"cd",  x"81",  x"fe",  x"67", -- 0D50
         x"cd",  x"89",  x"fe",  x"6f",  x"d1",  x"c1",  x"c0",  x"c5", -- 0D58
         x"0e",  x"01",  x"af",  x"cd",  x"83",  x"fe",  x"f5",  x"84", -- 0D60
         x"67",  x"f1",  x"85",  x"bf",  x"cd",  x"89",  x"fe",  x"6f", -- 0D68
         x"c1",  x"c0",  x"db",  x"88",  x"5f",  x"7d",  x"fe",  x"48", -- 0D70
         x"28",  x"6e",  x"fe",  x"41",  x"28",  x"06",  x"fe",  x"46", -- 0D78
         x"20",  x"0d",  x"3e",  x"a9",  x"d6",  x"2c",  x"6f",  x"7c", -- 0D80
         x"fe",  x"38",  x"c0",  x"7d",  x"c3",  x"38",  x"fe",  x"fe", -- 0D88
         x"40",  x"28",  x"6b",  x"d0",  x"d6",  x"39",  x"d8",  x"84", -- 0D90
         x"cb",  x"78",  x"28",  x"2d",  x"01",  x"90",  x"00",  x"26", -- 0D98
         x"05",  x"ed",  x"61",  x"0c",  x"ed",  x"60",  x"0d",  x"ed", -- 0DA0
         x"41",  x"cb",  x"7c",  x"c8",  x"3c",  x"fe",  x"0c",  x"38", -- 0DA8
         x"64",  x"28",  x"60",  x"fe",  x"0e",  x"38",  x"5e",  x"28", -- 0DB0
         x"5a",  x"fe",  x"0f",  x"28",  x"58",  x"d6",  x"2b",  x"38", -- 0DB8
         x"4e",  x"fe",  x"0d",  x"d0",  x"21",  x"33",  x"fb",  x"18", -- 0DC0
         x"55",  x"3d",  x"d6",  x"0a",  x"d8",  x"d6",  x"06",  x"c8", -- 0DC8
         x"30",  x"0d",  x"fe",  x"fa",  x"20",  x"02",  x"d6",  x"1f", -- 0DD0
         x"cb",  x"73",  x"c8",  x"d6",  x"80",  x"18",  x"38",  x"fe", -- 0DD8
         x"1b",  x"38",  x"34",  x"fe",  x"1e",  x"c0",  x"18",  x"2f", -- 0DE0
         x"7c",  x"fe",  x"0c",  x"38",  x"26",  x"28",  x"26",  x"fe", -- 0DE8
         x"0e",  x"38",  x"20",  x"28",  x"20",  x"d6",  x"2b",  x"38", -- 0DF0
         x"18",  x"21",  x"40",  x"fb",  x"18",  x"20",  x"78",  x"a9", -- 0DF8
         x"ba",  x"c0",  x"3e",  x"03",  x"a4",  x"7c",  x"20",  x"c2", -- 0E00
         x"b7",  x"20",  x"a2",  x"3e",  x"5f",  x"18",  x"08",  x"c6", -- 0E08
         x"20",  x"c6",  x"2b",  x"c6",  x"10",  x"c6",  x"20",  x"cb", -- 0E10
         x"73",  x"28",  x"1d",  x"21",  x"53",  x"fb",  x"06",  x"00", -- 0E18
         x"4f",  x"09",  x"7e",  x"fe",  x"5e",  x"28",  x"f0",  x"fe", -- 0E20
         x"5d",  x"28",  x"ec",  x"b7",  x"e1",  x"20",  x"0a",  x"3e", -- 0E28
         x"7f",  x"32",  x"24",  x"00",  x"3e",  x"0a",  x"18",  x"43", -- 0E30
         x"e1",  x"fe",  x"7e",  x"20",  x"0d",  x"7b",  x"ee",  x"40", -- 0E38
         x"d3",  x"88",  x"af",  x"32",  x"24",  x"00",  x"3e",  x"28", -- 0E40
         x"18",  x"31",  x"fe",  x"7d",  x"20",  x"0a",  x"3a",  x"26", -- 0E48
         x"00",  x"ee",  x"01",  x"32",  x"26",  x"00",  x"18",  x"ea", -- 0E50
         x"c1",  x"d1",  x"e1",  x"fe",  x"5d",  x"28",  x"06",  x"fe", -- 0E58
         x"60",  x"20",  x"03",  x"d6",  x"21",  x"3c",  x"b7",  x"c9", -- 0E60
         x"3e",  x"83",  x"d3",  x"93",  x"af",  x"d3",  x"90",  x"3e", -- 0E68
         x"25",  x"d3",  x"82",  x"3e",  x"96",  x"d3",  x"82",  x"af", -- 0E70
         x"32",  x"24",  x"00",  x"32",  x"23",  x"00",  x"af",  x"18", -- 0E78
         x"d7",  x"3e",  x"f7",  x"06",  x"08",  x"81",  x"cb",  x"3b", -- 0E80
         x"d8",  x"10",  x"fa",  x"c0",  x"81",  x"bf",  x"c9",  x"f3", -- 0E88
         x"db",  x"91",  x"2f",  x"57",  x"3e",  x"03",  x"d3",  x"93", -- 0E90
         x"3e",  x"fb",  x"d3",  x"90",  x"db",  x"91",  x"67",  x"3e", -- 0E98
         x"fe",  x"d3",  x"90",  x"db",  x"91",  x"6f",  x"3e",  x"cf", -- 0EA0
         x"d3",  x"92",  x"3e",  x"ff",  x"d3",  x"92",  x"3e",  x"cf", -- 0EA8
         x"d3",  x"93",  x"af",  x"d3",  x"93",  x"d3",  x"91",  x"db", -- 0EB0
         x"90",  x"2f",  x"5f",  x"3e",  x"80",  x"d3",  x"91",  x"db", -- 0EB8
         x"90",  x"2f",  x"32",  x"13",  x"00",  x"3e",  x"40",  x"d3", -- 0EC0
         x"91",  x"db",  x"90",  x"2f",  x"32",  x"14",  x"00",  x"cd", -- 0EC8
         x"15",  x"fb",  x"af",  x"d3",  x"90",  x"c9",  x"f3",  x"af", -- 0ED0
         x"32",  x"69",  x"00",  x"cd",  x"0a",  x"fb",  x"d3",  x"93", -- 0ED8
         x"cd",  x"0d",  x"ff",  x"cd",  x"31",  x"ff",  x"ed",  x"a1", -- 0EE0
         x"ea",  x"e3",  x"fe",  x"cd",  x"29",  x"ff",  x"3a",  x"6b", -- 0EE8
         x"00",  x"cd",  x"18",  x"ff",  x"2a",  x"1b",  x"00",  x"06", -- 0EF0
         x"80",  x"7e",  x"cd",  x"18",  x"ff",  x"3a",  x"69",  x"00", -- 0EF8
         x"86",  x"32",  x"69",  x"00",  x"23",  x"10",  x"f2",  x"cd", -- 0F00
         x"18",  x"ff",  x"7a",  x"18",  x"2b",  x"3e",  x"85",  x"d3", -- 0F08
         x"80",  x"3e",  x"40",  x"d3",  x"80",  x"fb",  x"57",  x"c9", -- 0F10
         x"c5",  x"4f",  x"06",  x"08",  x"cb",  x"09",  x"f5",  x"dc", -- 0F18
         x"31",  x"ff",  x"f1",  x"d4",  x"2d",  x"ff",  x"10",  x"f4", -- 0F20
         x"c1",  x"1e",  x"80",  x"18",  x"06",  x"1e",  x"20",  x"18", -- 0F28
         x"02",  x"1e",  x"40",  x"7a",  x"cd",  x"38",  x"ff",  x"7a", -- 0F30
         x"32",  x"6a",  x"00",  x"3a",  x"6a",  x"00",  x"b7",  x"20", -- 0F38
         x"fa",  x"53",  x"c9",  x"f5",  x"3e",  x"03",  x"d3",  x"80", -- 0F40
         x"3e",  x"85",  x"d3",  x"80",  x"3a",  x"6a",  x"00",  x"d3", -- 0F48
         x"80",  x"af",  x"32",  x"6a",  x"00",  x"f1",  x"fb",  x"ed", -- 0F50
         x"4d",  x"f3",  x"cd",  x"0a",  x"fb",  x"d3",  x"93",  x"d3", -- 0F58
         x"8a",  x"3e",  x"05",  x"d3",  x"80",  x"3e",  x"b0",  x"d3", -- 0F60
         x"80",  x"3e",  x"0f",  x"d3",  x"8a",  x"3e",  x"0a",  x"d3", -- 0F68
         x"8a",  x"3e",  x"e7",  x"d3",  x"8a",  x"fb",  x"06",  x"16", -- 0F70
         x"cd",  x"d1",  x"ff",  x"38",  x"f9",  x"fe",  x"90",  x"38", -- 0F78
         x"f5",  x"10",  x"f5",  x"06",  x"02",  x"af",  x"32",  x"69", -- 0F80
         x"00",  x"4f",  x"32",  x"6a",  x"00",  x"cd",  x"e0",  x"ff", -- 0F88
         x"fe",  x"52",  x"30",  x"f1",  x"10",  x"ef",  x"cd",  x"e8", -- 0F90
         x"ff",  x"d8",  x"32",  x"6b",  x"00",  x"06",  x"80",  x"2a", -- 0F98
         x"1b",  x"00",  x"cd",  x"e8",  x"ff",  x"d8",  x"77",  x"3a", -- 0FA0
         x"69",  x"00",  x"86",  x"32",  x"69",  x"00",  x"23",  x"10", -- 0FA8
         x"f1",  x"cd",  x"e8",  x"ff",  x"d8",  x"47",  x"3a",  x"69", -- 0FB0
         x"00",  x"b8",  x"c8",  x"37",  x"c9",  x"f5",  x"db",  x"80", -- 0FB8
         x"f5",  x"3e",  x"07",  x"d3",  x"80",  x"3e",  x"b0",  x"d3", -- 0FC0
         x"80",  x"f1",  x"32",  x"6a",  x"00",  x"f1",  x"fb",  x"ed", -- 0FC8
         x"4d",  x"af",  x"32",  x"6a",  x"00",  x"3a",  x"6a",  x"00", -- 0FD0
         x"b7",  x"28",  x"fa",  x"4f",  x"af",  x"32",  x"6a",  x"00", -- 0FD8
         x"3a",  x"6a",  x"00",  x"b7",  x"28",  x"fa",  x"81",  x"c9", -- 0FE0
         x"16",  x"08",  x"af",  x"5f",  x"cd",  x"d1",  x"ff",  x"3f", -- 0FE8
         x"30",  x"04",  x"fe",  x"90",  x"d8",  x"37",  x"cb",  x"1b", -- 0FF0
         x"15",  x"20",  x"f1",  x"cd",  x"d1",  x"ff",  x"7b",  x"c9"  -- 0FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
